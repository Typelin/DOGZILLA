MZP      ��  �       @    ��jr                             � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                                                                                                                                                                                                                                                                                        PE  L Ȅwh        � #  �        x      �    @                      �         @                      � L    � |   �  
                  �  	                                                                                  .text    �      z                    `.data      �   ,   �              @  �.tls        �     �              @  �.idata      �     �              @  @.edata      �     �              @  @.rsrc      �  
  �              @  @.reloc      �  
   �             @  P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �&@  �>@  �<@  0D@  ��G@  �W@  �Y@  |[@   @]@   �b@   tf@    i@   �i@   �@   �?@  �[@  _@   �b@   8i@       �fb:C++HOOK���@ �@ ���@ �����@ �D$�	�@ ����@ �=	�@ ud�=��@  t$�w  ���@ %   �t�Đ@ R�5  X3��   ���@ �=	�@ u ��H  R�T$���@ �!  Z��  �!  j �-V  YhL�@ �D$���@ �=	�@ t�=	�@ t��F  ���@  ����@ �=�aA  tP�	�@ P�D$P��aA �=��@  t�F  ���=	�@  u�Q  � !  �+H  ��   � ��U  3����@ á��@ �`� P��Sh�  ù�   �tQ�=��@  s
��   �������   Qj��u  P��u  �u
��   ����WVPP�5��@ �KH  �5��@ �TH  _^_ù�   �t�H  ���@ �� s���   �v���Ã=��@  r(�5��@ ��G  �tPj�]u  P�{u  �5��@ �H  �Ã=��@  t�����5��@ �G  Ã=��@  u
�G  ���@ �5��@ �G  ��t��������@ P�G  á�I@ ���U���ܸ0�@ �J  �UR�   Y�M�d�    ��]�U���ܸ@�@ S�]�\J  ��tS��  Y�U�d�    [��]Ð��o8  Ð��=L�@  t�L�@ �X8  Ð���=P�@  t�P�@ �����Ð��U���ܸ\�@ S�]��I  �M���t�t�@ ��EtS�j���Y�M�d�    [��]Ð�U��T�@ ]Ð�    0     s   @ D                   P@  H std::exception                  0     w   @ P                   �@  T std::bad_cast   �@                    U���ܸ��@ �I  f�E� �t�@ �M��E�d�    �E��]�     �@ std::exception * ���U���ܸ��@ S�]�H  ��t�M�j S�������EtS�&���Y�U�d�    [��]Ð�3�ÐSV�������@ �؅�tVj S�  ����^[Ðh̑@ ��r  ;��@ thՑ@ �2  YÐ�U��SVW�}�u��t�} t�} u3���   h�@ �Yr  �؅�u3���   h�@ S�Mr  �h'�@ S�@r  �U�hB�@ S�0r  �M�ha�@ S� r  �h|�@ S�r  �U�h��@ S�r  �M�����@ �? u��@ �E�8 u	�U��@ �M�9 u	�E� �@ �> t%�U�: t�M�9 t�? t�E�8 t�U�: u3���   _^[]�SV������@ �  ��u3��(  hڒ@ �bq  ���5��@ ��u3��  �����T$R�L$Qh��@ h��@ h��@ h��@ ������h�@ ���@ Q�q  ���@ h��@ ���@ P�
q  ���@ �=��@  t	�=��@  u1�C�1@ �C2@ �C 2@ �Ct2@ �C82@ �C   �   �r�=��@  t�=��@  t	�=��@  uh�@ �0  Y�{ u�{ thX�@ �|0  Y�Cd@ �Cx@ �C�@ �C�@ �C�@ �C   ���@ �   YZ^[ÐU��E��t���@ ]Ð�U��E��t���@ ]�3�]Ð�U��E��t���@ ]�3�]Ð�U��E�U��u��t&���@ ]����u
�����@ ��ȋ����@ ]�3�]Ð���@ ÐU��EP���@ Y]�U��EP���@ Y]�U��������u<���@ �1@ ���@ 2@ �ȓ@  2@ ���@ t2@ �ē@ 82@ ���@    �E���@ ]Ð�U��j����Y�EP���@ Y]�U��j����Y�EP���@ Y]�U��j�r���Y�EP�ȓ@ Y]�U��j�Z���Y�EP�UR���@ ��]Ð�Ð�����@    Ð�=��@  t�ē@ �3�Ð��tjPh�@ ��  ��Ð����@ �*)@ ;u6��,@ ;Hu,��.@ ;Pu"��1@ ;Hu�l@ ;Pu�p@ ;Hu3���   Ð���@ �T&@ ;t6�h&@ ;Ht,�|&@ ;Pt"��&@ ;Ht�l@ ;Pt�p@ ;Ht3���   Ð�S���&�=ғ@  uj �n  �˲3���  ��tj
�kn  �˲3���  ��u�[�S�=Г@  t3ۋ������@ ����C��7r�[�S���  jh   h�� j �?n  ��tM���@ � ��@ ���@ �P��Ё��� ��+Ӄ����   ��� +˃�����@ � �@ �[�[�3���@ 3�[Ð�=Г@  t
���@ �����SVW����  N����  ��jh  Vj �m  �؅�t.�{���s�������@ ���@ ���@ �C����@  ����_^[Ð�SVWU��������{����.�F�$�Fuh �  j V�Hm  ��t3��B����=�F�ރ��3���j�D$PS�(m  h �  j S�m  ��u�����D$;�v+���υ�u�$�*�$�M���@  �ǃ� ]_^[Ð�SVW����U������ڋ �������;���   �����;�v�����׃����Љ$j�D$P�L$Q�l  �|$   un�d$  ����+֋D$;�sZ��+΁�   I��  ����;�s��jh    V�D$P�<l  ��t+jh   V�T$R�&l  ��t�ǃ��Xp���p���|����  ����tm��,
 v�ƃ��X�׃��B�ȋ֋��`  ���.  �A��;�r
�����_�1����  ����t"��,
 v�ǃ��X�͋֋��J  ����  �ƃ� ]_^[Ð���ȋу�����ыȃ�������u3��Ð���@ ��t� �@ ;�r�ȁ��� ; �@ s���Á��� t� �@ �3�Ð�S�؃� V��;Bu�Z;Zv���ރ�������B+؉^[Ë�ZK�^[�3�Ð3�ÐSVW��h�  j S�  ��3ҋù�@ �1�0�1����p�x }3��pB���� ��7|������=Г@  t
���@ ������5��@ �l��x  �� ��������tT�Ѓ����u?�ʃ����t&����@ ������)�x  ��L;�HL���p  ���t  ������u��v����@ u����@  3Ҹ�@ �  B�� ��7|��
������@ ��P�����|  ��  �H��  �@=��@ u����@  _^[Ð��SVW����h   j V��  ���=Г@  t
���@ ��������@ �����3ۍ�C��r�R����@ u����@  �r������@ �#�J�����3���<C�>����;�r�R����@ uՋ����@  ��3ۀ> u.j�T$R����Q�	i  �|$   u���|$    u�CF��   rÃ�_^[Ð�SVW��ԉ$�t$j(j V��  ���1����=Г@  t
���@ ������=��@ �   �   �F   �F  ��������ta�Ѓ���ʃ����uD��t3����@ �������@ �X����+ʃ�N�KN +�V���N�F �N������u������@ �t�����@ F���@  3Ҹ�@ �  B�� ��7|���������@ ��P���V�HN+�V �@=��@ u����@  �~~~�~�$V���
   �^�$��,_^[Ð���u3�Ã�� �u� �P������èu������èu�������3��SVW�����u3��  �ȋу����u/��X�����;�r����@;�w
�   ��   3���   ��   ��um�ڋу���ƃ�Ӄ�;�s�����tH����;�r?�   �   �3���;�w�   �   ���,  |	�   �z�=�  r�   �j3��f�d��u]�ڃ������;�s<������j�T$RP�tf  �|$   u�d$  ��+�;|$s�   �3�����;�r�   �3���3���_^[Ð��S�>e  ��3�������������@ �   +؈���@ @��|�[Ð��SV�����h��@ j j�e  �؅�u3�^[�j j j jS�le  �0P�e  S�d  ��^[Ð���S�����u[�=��@  uL���@ ;��@ u&���@ ;��@ u������t�����   �3���h   he�@ h(�@ j �oe  3�ø   �3�ÐS�������uS�=��@  uJ�<�����u=h��@ jj jj j��d  j j j ��jS���@ �d  � ԓ@ P��d  �   [�3�[�3�[Ð��VWU��@ 3�3��=��@  t�����Du-�����t��y������������@ ;�v�
@B;�w���G��7r�]_^à��@ Ð�Q�$�$:��@ t�$���@ ����ZÐSVW�=ӓ@  �f  �ӓ@ �<�����t
�ԓ@ �����3��8�@ �; u��'@ �Ƌ���3������@ �C����@ �S�K��C�   �K�����@�   % �����0=0  s�0  �  ����v�   �Ȳ������S�f0f�C��{�����I���   �� �����0��0s  s�0s  ��0�  v�0�  ���� 3����S���f��� f�� �f��0f�S�F�� ��7�����h������@ ��@ ���@ ��@ 3���������@ � �@F��   |����@ ��@ ���@ ��@ j �Hb  ;��@ u������>���_^[Ð�SV���@ WU���@ �F��@ ��hh �  j P��b  ��;�u�3ҍC����ˉ����ˉH�3��@�   �H�B�� ��7|؉6�v3ҋ�������@ � �@B��   |�G��Xh �  j P�Xb  ��;�u�?�]_^[À=ӓ@  t6�ӓ@  ���@ ��tP�a  3҉��@ �4���������u
��@ �����S����������  [Ð��S���������7  [Ð��SV����q����֋��  ^[ÐS���\������  [Ð���K���Ð���Ë�
�H�@�J�BË�
�H�J�H�J�H�@�J�BË�
�H�J�H�J�H�J�H�J�H�@�J�B��(�h�h�h�H �J �z�z�z�:��(�h�h�h�h �H(�J(�z �z�z�z�:��(�h�h�h�h �h(�H0�J0�z(�z �z�z�z�:��(�h�h�h�h �h(�h0�H8�J8�z0�z(�z �z�z�z�:��(�h�h�h�h �h(�h0�h8�H@�J@�z8�z0�z(�z �z�z�z�:Ã�����y�,�l�|
�<
��x��,�<
�D�D
Ã������,�<
��x���
ËH�;ʉ�JtÐ�錽@ �����ָ������!��@ u���������!�@ Á�0  �����  �#с��  �Ռ�@ �Q;щ�P��AtÐ��錽@ �����ָ   ��	��@ �   ����	�@ Ã=�@  uÐ�� �@ �@�u%�H���@ +J�H��T���0  �g���Ð������#P���0  r����� �@ �����#P���@ +���ÍP��=,
  S�Г@ �H  ������@ ���@ uV�S�B�����;�t�B#H��J�P�t(� [Ð���S�K�;Cwv�B�K� �P�[Ð���J�Y�K� [Ð��   ��#t��� �   ��#t��� �   ��#t���@�=ғ@  u�j �L^  �   ��#�_���j
�6^  �VW�=Г@  t9�   ��%��@ t*�=ғ@  u�j �^  �   ��%��@ t	j
��]  ���s#5�@ tp�ƍ4�    ���@ �ɍ��<͌�@ �w�V�W�:;�u�������!��@ u��@ �����#~���`
 rl���{+׍>�J�H��T������U�K�=�@ ;�r&�5 �@ �K��0  ;�r��+�)=�@ �5 �@ �!�C�����������u���@ �_^[Àd>���O�N�3����@ ��F�F   �s�F �K��S�+��{� �p�_^[Ð�   ��%��@ tK�=ғ@  u�j ��\  �   ��%��@ t*j
�\  �ǐ��=,
 �  ���   �� �����0��u��������������������#��@ t�������^�����������#�@ t�Ћ��@ �ȋ�����5���@ +�r� �@ +ã �@ ��@ ���X������������@  [�VW�<͌�@ �w�F�G�8;�u�������!��@ u��@ �����#~���+�t��J�H��T���0  r����������d>���K�N����@  ��_^[�[�������3�ËP�����S�Г@ ��   �ۋua�j�Bt,���J�@�A�t3��[Ð�K�Z�J�Q�S� 3�[Ð���t�B�J�H�A3�9Su�C��R��Г@ �   �   ��#t��=ғ@  u�QRj ��Z  ZY�   ��#�o���QRj
��Z  ZY�Ð���   ��%��@ tB�=ғ@  u�j �Z  �   ��%��@ t!j
�Z  �ǐ������   ����ۋ�V��u��D�   �L�u5���L��F�u@���� tP�C�F��\��Ƌ��n������@  3�^[Ð����ف�0  r�����뻐�N�+�ف�0  r��������먁=�@ �� u,����V�P����@  h �  j V�Z  ���^[Ð������ �N����C�   ��@ �� � �@ ���@  3�^[Ð�[���H��������ËH���SV����   ��K��;�r7��@   ;�r^[Ð�ڋ��O�����t�ˋЋ؋�������������^[Ð��L	 W��3�+ʃ��#��������t$��,
 v�x��K���Ћ����S���w�����_^[Ð���k  �ك��W�<����;�U�  �,;�r]_^[Ð����,  s���  ��   �,  ;�vۍ��   �� �����0��+̀=Г@  tF�   ��%��@ t/�=ғ@  u�Qj �hX  Y�   ��%��@ tQj
�PX  Y�Ð�   #^�݉^��ًW���u	���W����ǃ������0  r�����_��C�D.���0  r
�.���'������@  ��]_^[Ë����������t��ЋƋ��������G�����]_^[ËG����   ����,;���   �=Г@  t_�   ��%��@ t3�=ғ@  u�QRj �W  ZY�   ��%��@ tQRj
�eW  ZY뿐�   #^��G���~   ����,;�wt=0  r��QR�"���ZY�����3�+��#Ǎ��   % �����0�U+�w�$.�������T.��z�|����0  r������n����@  ��]_^[Ð����@  �����3�+��#���R����Z��tс�,
 v�P���ЋƋ��6�����������]_^[Ð^[�������3��S�X�����^�����ɍف�,
 s�������x��
����[Ð�U��E��t��@ ]Ð�U��E��u3�]���@ ]Ð�U��E��u3�]���@ ]Ð������Ð�U��S�]��t�U��������t��[]�3�[]ÐU��E�]���]Ð��U��U�E��u��t��@ 3�]Å�u
����@ ]���@ ]Ð��Ð��Ð��Ð��U��3ҋE�B��f�8 u���]ËT$�D$�L$�   �D$Ð�;�t5�� �|   ���$�@3@ �,�(��~�h��~�h�z�z�:�<
Ð�3@ �3@ �3@ �3@ �3@ �3@ �3@ �3@ �3@ R�(�D��L��(Q�ك���LZ�,�<
��|��:Z�:�~.;�w�+�;
vȃ�Q�,�(ʃ��+��,�<
���Y�:�<
���
��f�
�f��@f�
�BË�
Ë�@�
�BËf�@�
f�BË�@�
�B��(�:ËT$�D$�L$������D$Ð�� ��|?f�f�Hf�Hf�H��� ��T�ȃ���+�������T��|�����Ð����~P�L�����ڍU�4@ �␐f�Hf�Hf�Hf�Hf�Hf�Hf�Hf�Hf�Hf�H
f�Hf�Hf�Hf�Hf��ÊL$�T$�D$�T����D$��萋T$�L$3�8t8Bt8Bt8Bt��8��BBB����t(�A�B��t�A�B��t�A�B��t
�����Ґ��D$Ð���D$�u-����ʁ�� ��t���#�t��u(��u%��  � u����@��t�@��t�@��tH$��HHH�L$H+�Ð��D$�T$�L$IxjS��3�8t8Ct8Ct8Ct����CCC����t<Ix4�B�C��t/Ix&�B�C��t"Ix�B�C��tIx
�����Ɛ�CCCC3��[�D$Ð�U��S�];<�@ r3�[]Ë�l�@ R�Q  ������[]Ð��U��EP�fQ  ������]ÐU��SVW�];<�@ r
j��  Y�d�E��rt	Ht�3���   ��   �
j�  Y�9S��  Y�$�@�@ ����Wj �EP��l�@ R�Q  ��@u��  S�D  Y��_^[]�U�������SVW�}�E;<�@ rj��[  Y�  �UB��s3���   �UR�h  Y�M��A�@ tjj �EP�!������U��A�@ @u�MQW�EP��   �����   ��3��E�3҉U��{��������F<
u�E��C�
C��C��������+ʁ��  }	��+�;Mr΍�������+Ѝ�����RQ�EP�b   ��������+�;�t���u���� �]�+]���E���+�;E�x����]�+]��EP�  Y��_^[��]Ð�U��E��t�  3�]Ð��U��Q�E;<�@ rj�  YY]�j �U�R�MQ�UR��l�@ P�7P  Ht�c  Y]ËE�Y]Ð�U��EP�UR�MQ�\�����]Ð��U��SVW�]�}�u�Ct
�CP�~���Yf�c��3҉S�K�K��}t>��v:��@ �A@ ��uW�<���Y����tf�K������3�s�{�}uf�K3�_^[]Ð��U��SV�]��u	�   3��v:[t����lS�o  �{ Y|"�Cu�S;u3ɉK�K;u�C�3��4�ssF)sV�C�P�SR�k�����;�t�Cu
f�K����3�S��  Y��^[]ÐU��E���@����@ ]ø��@ Ð�SVWU�  3�=<�@ ��������7�C��}-�s�F)sV�C�P�SR�������;�t�Cuf�KE���σ����u��y  ��]_^[Ð�U��E��@ ]Ð��U��E��t� ���@ ]Ð�4�@ P�"  YÐ���8�@ ��tP�����Y3҉8�@ ��@    Ð�4�@ P�q"  YÐ��U��SV�]�8�@ ��t�<� ui�����=8�@  u6�5<�@ ��V�\���Y�8�@ ��uh�@ �4"  YVj �8�@ R��������8�@ �<� uh1�@ �����R�|!  ���p����8�@ ��P��!  Y^[]�U��SV�u3ۃ=8�@  uh�   hM�@ hF�@ ��	  ���=�@  t�8�@ ��R�"  YHu�   �8�@ ��R�!  Y��t�����^[]Ð�U��3��@�@ �	�: t@��;<�@ |�;<�@ u���]ËU��@�@ �M��l�@ ]�U��E�M���u3��@�@ �@��;<�@ }�: u�<�@ ;�v;�w���]Ë�@�@ ��t
�<�@�@  t���]É�@�@ �M��l�@ ]�U��E;<�@ s	3҉�@�@ ]Ð��U�����<�@ ��V�u��<�@ t�: uH�����u��u��u3��b�������X�3ɉM����E�@�@ ;E�~.��U����t�� �ƀu�ɀ�� t��@�F�E��E�;E����Phl�@ V� �����3�^YY]Ð�SVW�ĴhW�@ h4�@ �  ���<�@ P�KK  ��;<�@ s�<�@ ���@ <@ 3҉T$�L$Q�J  �D$:�t$<����   ��$���$����;���   �D$   3ۿ@�@ ;$}<�F3��� t   ��@t    �t @  � �  ���ȉC��;$|ċ$��@�@ �3�C���;<�@ r��$��QVhl�@ �8������|$ uej��J  �l�@ j���I  �p�@ j���I  �t�@ 3۾@�@ S� ���Y��u	�=��@  t�    �=��@  t�   ��&����C����~ƃ�L_^[Ð�O  ��Ð��U��S�]��|��*  v�   ��������t�@ �����;h�@ }������ �����  ����[]�S�I  �؁���  ��%��  P����Y��[���H  %��  P����YÐ�Sh8�@ h<�@ �  ��������3��Q��@���[و����r�   �Q^��������[وZ@��;<�@ r�j �_����@Y��A�@  uj �I���Yf�`��h   j �6����@Yt�   �3�Rj j ����YP������j�����@Y��A�@  uj�����Yf�`��h   j������@Yt�   �3�Qj j�����YP������[��   j �����@Yt;j ����YP����Yj ����Y�@P����Yj ����Y3҉Pj �t���Y3ɉHj�g����@Yt;j�Y���YP�����Yj�J���Y�@P�����Yj�8���Y3҉Pj�+���Y3ɉH�   Ð���<�@ P�Y  YÐ���<�@ P�Y  YÐ��U��SV����P�EZ+¹   ����ء@�@ ��t�<� ui�����=@�@  u6�5<�@ ��V�1���Y�@�@ ��uhT�@ �	  YVj �@�@ R�������@�@ �<� uhq�@ �����R�Q  ���]����@�@ ��P�  Y^[]Ð�@�@ ��tP�����Y3҉@�@ �4�@    ÐU��SVW3��}�4����؃=@�@  uh'  h��@ h��@ �q  ���=4�@  t$��+ù   ����@�@ ��P�  YHu�   ��+ù   ����@�@ ��P�  Y��t�X���_^[]Ð��SV����3���������CtS�����YF��;5<�@ r��h���^[ÐU��e��}����E���]ÐU��e���}��M��E���U#���#��f�E��m����@ ��]Ð��h�  �5��@ ���������Ð��U����SVW�}�u�]��|M��$H��}�} t�-C�ލM܋�3����A��3�������t��I�<
}��0�C�E��C�U�;�u�� �E_^[��]Ð��U��jaj j
�EP�UR�v�����]ÐU����SV�u���u	�D  ������u	�YD  ������u�Ԩ@ �0��t!�E�PV�AD  ��uh �@ �9  Y�����   3��D�@ � @B=  |����   �}���   �M��3ۊ؋Í�E�@ ��@B3ۊY;�~�����t�y uՁ��  uj�@   ���@ �
@B��~~���   ���@ �
@B=�   ~�3����@ ��E�@ ��
@B3Ɋ��@ ;�~�3����@ ��E�@ ��
@B3Ɋ��@ ;�~�5H�@ �3��H�@ 3�^[��]Ð��H�@ Ð��7C  P����YÐ��U��SV�M�E3�3ۊ��E�@ t'�x u@��u-���)� 3ۊ���p�;�u��@�
3ۊ;�u�Њ@��u���^[]�U��QSVW�]� �E�E��S�]���Y�}+�O��~WVS�������E��E��p���u�_^[Y]Ð��U��j h_�@ �EPhW�@ �URhD�@ h�   hL�@ ������ hL�@ �����Y��L�@ P�MQ������hL�@ �B  Y�P  ]Ð����T�MB  �D$P�T$R�L$Q�D$P�T$R�L$Q�D$Phh�@ hL�@ ��B  ��$�L�@ ��Ð�U��QSVW�}j h�   jj j h   ��EP�A  �؅�u�7�~������E�j PV�@���YPVS�B  j �U�RW�+���YPWS�zB  S�TA  _^[Y]Ð�SV�A  ���n  ��V���B  ��^[Ð�U��E�    3�]� ��Q3��$�A  ��f%�����ƀu�    ZË�RhF@ � A  P�B  �<$ t�    ��   Z�U���|����=��@  SV�u��   �=��@  ��   �=��@  tch�   ��|���Pj ��@  j\��|���R�v������؅�uj:��|���R�_������؅�u��|����C�8���  PSVj �oA  �   j��@  �؍E�j Pjh��@ S�@A  j �U�RV�����YPVS�+A  j �M�Qjh��@ S�A  �;�=��@  t�=��@ �t)V���@ Y���@ ��t�=��@ �t�8 t
VP������^[��]ÐU��EP�����Y]ÐU��EP�����Yj�  Y]Ð��@ �h�@ ÐU���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������]Ð��U���ظ��@ SVW�  3҉U�f�E� �M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�i���f�E�  ��x�   �M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�M�Q�E�P�U�R�������x�M�d�    _^[��]Ð�U�존�@ �U���@ ]ÐhЪ@ �Z���Yj�  Y�U���ܸ��@ SVW�  f�E� �=��@  t�<  ��tj j j h  @�<  f�E�  ��}�  @�����������}Ћuԋ]�]Ðj�a
  Y����Ð�U����3�SV�]�M�E�����E����;U�~�8 u�;E�tR�U��E�@�ӉU����@��;}�: t�;u	�E���(��Ëu���T��u��V3҉�3҉T��E��E��^[YY]�U��SV�]�u�  �;   u�  �   ���M�L���E����t  3�^[]Ð�U��hl!A hl�@ �EP�UR������]ÐU��hpaA hp!A �EP�UR������]ÐU��QSVW�}�  �E��U��u�N�E����|(���t;�t���u3҉�S�M�	;M�uN�����}؅�}ƋEP�UR��������
  _^[Y]�U��hl!A hl�@ �EP�~�����]ÐU��hpaA hp!A �EP�b�����]ÐÐ��U��S�]�h
  ��u�EP����Y�!
  ��@ �} u��u���@ ���@ �D
  �UR�	  Y�5
  []Ð�U�졟�@ P�URj j ������]ÐU�졟�@ P�URj j�z�����]ÐU�졟�@ P�URj j�^�����]ÐU�졟�@ P�*���Y�UR�����Y]Ð���@ Pj jj �+�����Ð�����@ Pj jj������Ð��U��j �EP�U��]Ð��U��j �EP�U��]Ð��U����SVW�]��u��E�j �UR�U������< t�<	t��:"u�����<"t��u��:"u�����< t<	t��u�R�6���Y@P�
���Y��taA ����   h �@ ����Y�   3����� < t�<	t��: ��   ��M��D<"u%��
SV�  ����<"t��u��:"u����<*t<?u�   SV��   ���� < t<	t��u��� ���t�MQ�M�Q�H�@ ���j �E�P�U����: t���9 �J����   _^[��]átaA ��tP�)���Y3҉taA Ð��U��SV�]�E�3��BA�9\t��9"u7�ʃ����
�0�\� �������u��t ��"� ���	��\� ��ʃ����u�^[]Ð��U��S�E�U��9\uPR������[]Ë3ۊ��E�@ t�y t
�	��� ����	�� �[]�U����SVW�]��u��E�j �UR�U�����f�f�� t�f��	t�f�:"u(����f�f��"tf��u�f�:"u����f�f�� tf��	tf��u�R����Y���P�����Y��xaA ����   h$�@ �j���Y��   3����f� f�� t�f��	t�f�: ��   ��M��Rf��"u,��
SV�3  ���f�f��"tf��u�f�:"u%�� �f�f��*tf��?u�   SV��   ���f� f�� tf��	tf��u��f�  ���t�MQ�M�Q�L�@ ���j �E�P�U���f�: t��f�9 �)����   _^[��]Ð�xaA ��tP�����Y3҉xaA Ð��U��SV�]�E�3��B��f�9\t�f�9"uA�ʃ�����0f�\ � �������u��t'�f�" � ����f�\ � ��ʃ����u�^[]ÐU��S�E�U�f�9\u(PR�w�����[]���f�y t��f�	f�� ���f�	f�� �[]Ð��U��3��|�@ �M;
t@����
|���]ÐU����SVW�]�]��E�E�3҉U��9  ����t�F(��u
�   �  3�����  �B��   ��  ���   ��  ���   J��   �   ��  ���   ��qt3��   ��o��?����   �$��S@ �S@ 'T@ �S@ :T@ �T@ dT@ �   �E��   �   �   �   �E��   �   �   �   �E��   �   �   �   �E��   �   �n�   �E��   �I   �[�E�   �   �M�E�   �   �?�E�   �   �1�E�   �   �#�E�   �   ��E�   �   ��   �y�4���u3��m��u�   �b3҃���t
��t��u8�;���h?  ���@ Q�>������M�Q�E�P��|�@ R�֋u����!~ ��E�Pj ��|�@ R�փ��E�_^[��]Ð��U��} u�   ��   P��   Y�   ]� ���U��SVW�=P�@  �]u���A  S@ jhU@ �2  �P�@ S����Y��@u�|����    ����c��t��u�T�@ �I��  ����u����B�_(��u2j(�2���Y�؅�u�6����    ����3ҋ�3�B�����
|�_(���U��_^[]ÐU��SVW�]��t��u�T�@ ��e  ����t�~(��u�   �^S�����Y��@u�   �K����tA��u'�����r5��t0��t�	�'������ j�V���Y�3҉�3Ҋ���@ j RS�Ѓ�3�_^[]Ð�U��EP�`  Y]� ���U��EP�0  ]Ð�U����SVW�E�8 ��   �} t�E������E�������   ��E�   �E�   3���;u���   3��E��U�J�M��f�}�} �t�x��8�} t�P��P�U��} u��;]�s/��:Cu�S��;]�r���]����;�w��:Cu�S��;�v��E��E��U�
;M��u�;u��t���_^[��]Ð��=��@  u(���@    jh�aA ������jh�aA �������Ð���aA P��  YÐ����aA P��  YÐ��h��@ h�aA �]  ��ÐU��   ]Ð�U����SVW�]�u�}���E�   �u�u1��aA ��aA ��u"�K/  ��aA �VDR����Yj �M�Q�]������MQSW�FP��   ����u4��aA u,W����Yj�U�R�+�������aA ��tP��.  3҉�aA ��_^[YY]�U��� ����@   SVW�� ����E�ԫ@ ��=Ы@  tH3��� ����Ы@ h   R��aA Q�.  �� ���QSh֬@ �� ���P�p/  ���� ���R�]���Y�   _^[��]� ��U��E� dg�  ]ÐU����S�E��aA PQ�E��X@ �U���dg�  �d�    YX�Ы@    �MQ�URP�U���Ы@    �E�P����Y��[YY]� ��U��EP�UR�MQ�����]� Ð��Ð��迸����   �賸����    �S��P���3��D$�   �D$P��-  �|$,u�   j�D$P�T$R�R.  �o���\$��    �İ   [Ð�.  Ð�U��EP�.  ]� U��EP��-  ]� U��EP�UR��-  ]� U��]� �U��]� �3�ÐS������   ��u�   ��������   ��[Ð�S��aA P�  Y��aA ��t
���aA �j`�$���Y�؅�tj`j S��������tT�CH   3�3ɉSL�KX3�3��K,�C\�{P u�P�@ R�߼��Y�CP��uS����Y3���P�@ Pj �SPR�f�������aA Q�  Y��[Ð��U��S�]��aA P�^  Y��aA ���aA ��aA Q�S  Y[]Ð��h$�@ h�aA ��   ��ÐSV��aA ������   ����   S����Y�   �؋C8��tP�7���Y�C<��tP�)���Y�C��tP����Y�C4��tP����Y�CD��tP�����Y�C0��tP����Y�C@��tP����Y�CP��tP�ջ��Y�C(��tP�ǻ��Y��P輻��Y�����i���^[�U��Sh�aA ��*  �=��A 2  |
�EP�e   Y���A ���R���aA R�R+  ���A �]���I���aA �h�aA ���A �C+  []Ð�U��EP�*  ]Ð�U��EP�"+  ]Ð�U��İVW�@�@ �}��ǹ   󥤋UR�M�Q�������E�P����Y_^��]Ð�U��EP��*  ]Ð�U��EP�*  ]Ð�U��E�@@]�h�aA �*  ���A    Ð��S��X�C�D$�C�C�]@ f�C  f�C  �C    dg�  �dg�  [�dg�  �**BCCxh1���5T�@ SWVUP�p�p�p�p��#  ��]^_[���U����SVW�}�Guh  h�@ hϭ@ ��������E�@uh  h�@ h�@ ��������U�Buh  h9�@ h�@ �������M�Y]�3��tg�Cu\�} t�C����t3���   �U�VW��  ����t�}� t
�   �   �Ft�u��uWV�3�������t�   �u��듋U�Z]�3��t^�} t�C����t3���   �U�VW�p  ����t�}� t�   �(�Ft�u��uWV���������t�   ����3�_^[YY]�U����SV�X�@ �'���3�����A ��t��t�X��t
jP� ����Å�u�F��   |ыU�d�    ^[��]�U��VW�M�u�}3�3�;�~:uB@;����_^]�U��V�M�u�U3�;�~
:t@;�����^]�U����3�3�3�SVW�E��U�M��} t	�E�@uhc  h��@ h��@ ��������} t	�U�Buhd  h��@ hˮ@ ��������} t �M�Auhe  h2�@ h�@ �������} tB�u�u��  ����thi  hg�@ h=�@ �n������u�u��  ����t3��  �} t�u�u�  ����tho  h��@ hr�@ �&������U�Bu3��Q  3҉U��M�Y]�;���
  �C��   �}$ t�C����t3���   �U�u�E(s�E��Ct�6�}�W�u�  ����u?�G��   �u��u��u �u�u�u�uWV�b�����$����   ���E ��U��X�u�} t;uuj���   �} t>�} uh�  hï@ h��@ �;�����j j �u j j �u�uWV�������$��u��}� t;u�u�U�	U���E��u�M�M���������}� u�E��E�X]������E �U���}�t3ɉM�E�_^[��]�U��QSVW�}�u�? uh&  h��@ h��@ ���������u3��i�V�U��} t�M��	�M��uS��   ����t�E���   �7�Ct,�CÅ�t"�U�R�uj P�|�������t�M��   �����_^[Y]�h��A �o���Y���@ ���A h��A �Z���Y�đ@ ���A �j h��A �Q�����j h��A �B�����Ð�U��S�]��u�d�@ []�f�{ ujhx�@ hm�@ �������C�[]ÐU��SVW�u�]��uh�   h��@ h��@ �p�������uh�   h��@ h��@ �U�����;�u
�   �   f�Sf;Vu�;t3��rf�SfV�t3��a�{�f�{ uh�   h��@ h��@ ��������^�f�~ uh�   hĭ@ h��@ ���������CG;�t3��	��u�   _^[]ÐU��QSVW�E�u�];�u
�   ��   �{�V�U��M�#���th��   �e�   ;}�tF��u>�ǋU���   %   ;�t*�E�%   ��#���t3��   ��   �M�   ;}�t3��~�   �[�v�u����U�#���t(�K;Nt��u�KNt3��L�   �[�v�C���VS�P�������t�   �'��   t�E�t�Ctj�uVS�������3�_^[Y]Ð    0     w   @ P                   f@  T std::bad_typeid �@                    U��SV�u�]�} u�E�`�CÍURVj P�l�������t�E�A�CÍURVjP�M�������t�E�"�
�@ ��th�  h{�@ hA�@ �������3�^[]Ð�U���ܸ��@ S�]�8�����tj S�$������EtS譬��Y�U�d�    [��]Ð�=��@  u
���@  @ �=��@  u
���@ 8@ ÐhT�@ j �"!  P�(!  ���A �=��A  u
���A �@ ÐU���ܸ��@ SVW�����̫����   ����A �:u�5��@ jj��   ��j �����Y���@ f�E� ��f�E�  ��  ����_^[��]Ð��s�����   ����A �8u�5��@ jj�   �����@ ���L���Ð��U����S�]��������t���u�U�R�+   Y�]�h�   S������   P�H����������[YY]Ð��U��S�]������$   �Ȱ@ �Isr��C��@ []ÐU��   ]Ð�U��S�EP�E@@Pj h����,   []Ð��U��SVW�}�u�]�;���u3���   �=���t=���u�Ƌ��  �|����;�  �u�=̓@  th��@ �e���Y�=��A  t�URWVS���A ����u3��m�=��A  t�URWVS���A ����u3��L�=��A  t1���A ���t��u�=���r=���vWSVjj�������;  @u�K����   _^[]ÐU��E3҉�@�g@ P�u   Y]Ð�U��EP�y   Y]ÐU�졜�A �U���A ]Ð���A �g@ Ð���A �g@ ���A �g@ Ð����aA ��tP����YÐ����aA ��tP�y���YÐ��U��Edg�  �dg�  ]�U��Edg�  ;�u	� dg�  ]Ã��t�9t�	�� ����n  �������SVWj Rh�i@ P�U  _^[�U���]Å�t
�   ��Q�Ð��h��@ j �  P��  ���A �=��A  u
���A �@ �U��S�]S�ح��Y��u5���   w�^�����   t�X����K�����   �?�����   []�[]�U��S�]�'���;�   u������   �[]�S肭��Y[]�U��QSVW�u�}�uj VW��������t
�   �   �W�U��^�� tF�uj�vW�b�������t�   �j�v�^��u3��Z�uj VW�8�������t�   �@��t9�Et�   �.�E�u3��$��@t��u�E�u��u�E�u�   �3�_^[Y]�U��SVW�]�}���uu�� th�  h��@ hȲ@ �o������Àth�  h�@ h�@ �S�������td��KtKtKt"��t(�/Wj V�U���   j WV�U�   ��3ҋ��U�Wj V�U�v�$�@ ��tmh  h3�@ h*�@ ��������T��KtKtKt��t�!WV�U���7VW�U�0�׋��U�'WV�U� �:�@ ��th9  hI�@ h@�@ ������_^[]�U��U3���t
�@�
B��u�]�U��SVW�} �ut�   �3��Et�ˀ   ���A �8u#�u�t���Y��W����YPW�ujj �������ƀ   th{  hi�@ hP�@ �	�������NtNtNt��t!�(S�u�U���<S�u�U�3�ӋE�U�)S�u�U� �p�@ ��th�  h�@ hv�@ ������_^[]�U��S�]�Àth�  h��@ h��@ ��������KtKtKt��t�%�u�UY[]��u�U[]ËE�U[]��u�U[]ú��@ ��th�  h��@ h��@ �.�����[]�U�����б@ SVW�u0�����]��tf�F  褤����   蘤����t�S��3҉�   �����M ��   �q����U$��   �]��{��   �3t�C�3���0   �E�t	�U؋J�M؍NRQ����Y�EЋE�3҉�MЉY�EЋU�P�MЉq�E�f�x�U�f�E�f�B�UЋM؉J�MЋE�A�U�3��B(�U�3ɉJ,�M��AQj@ �EЋU �P4�MЋE$�A8�UЋE�B �UЋM�J$�M��AE �E��@DV�u�UЃ�RR����������A �9t
���A �8ufS�����U4Y���r�M4�q�E4�p�U4�r�M4�q�E4�p�U4�2�MЀyD t�EЃ�R��UЋB@PS�����YPS�U(��Rjj�\�����4�E�te�} uh)  hĳ@ h��@ �Q��������A �M�f�E� �u�u�u�EЃ�RP����f�E�  ��������f�E� ��  �Ủ��A 襢����   �M��M��E(�EċUЉU�Qjjh����  �E�d�    _^[��]�U���ܸ�@ SVW�]�,�����uh  hԳ@ h˳@ ������f�E� j�uSj �u�u�
���f�E�  ����0���f�E� �%  �U�d�    _^[��]�U��SV�]�{D t.�Ct$�C�5��A �SR�H,Q�p(PR�[������5��A �CD �{E tB�s<��uhZ  h�@ h۳@ ��������Ft�Ft�F,P�v(V�s@�������CE ^[]�U����SVW�]�C(;Eth�  hI�@ h-�@ �������S,;Uth�  hl�@ hP�@ �������{E th�  h��@ hs�@ �h������M�A�C<���U  �U�B��H  �M���A���KR�U�M��CE�U�
M�K@�F�>�E��0t
�v�V�U��t �CtWj �s@�����E�   ���  �E���   �0��   � t&�Cth�  h��@ h��@ �������E�   �@�uh�  h˴@ h��@ �������Cuh�  h�@ hҴ@ �t������M��	�M�V�s���������u'�E��E�V�s�u���������E��U�;U�t�E�   W�M�Q�s@��������   �C��   �C;Cth  h�@ h��@ �������V�s�W�������uV�s�u��������E��E�   �FtC�U�z uh7  h1�@ h�@ �������M�q�E�p�u��s@������E�   ���YW�u��s@�b������H� tW�U�R�s@�L����E�   ���+;{th_  hO�@ h8�@ �;�����W�u��s@�������}� u$�E�t�Ft�N,Q�v(V�u��<������CD _^[��]�U����3�SVW�E�U�J�M��E��U+P�U��M�Y�+  �ËU��M�<���U��f�y����r����   tSJ��   ��   ��   �U��M�D���A f�A SUVW�{   �{   �M����A �>���_^][�uf�F  �   ������   �E���F(;Eu;^0u��u��U��2��u��t�M�;1th 	  hr�@ hV�@ ���������U��V����YV�VY�G�M�����M���u��uU�RP�Z  ���E�� �y�@ ��thX	  h��@ h��@ �������߅�t	;]�����_^[��]�U��SV�u�]���*�C��u���&j �vP�v�v���������t���
���; u�3�^[]�U���ܸ|�@ SVW�}�u�]�����Cuh�  hR�@ h*�@ �������{( uh�  hv�@ hY�@ �������f�E� f�E� ��t�U�J;K s*��u�M�A;C$s��uh�  h�@ h}�@ ��������   u��t�S ��S$�E)PV�K,Q�s(WS�u����f�E� ����-���f�E�  �"
  f�E�  �����f�E� �

  �E�d�    _^[��]�U��SVW�u�]�}�-�Cǃ} t� ��Bt�u$�u j V�uRP�   ��3���;]s�_^[]�U����SVW�u�E�@uhE  h?�@ h�@ ��������} t�U�Z ��E�X$��t;�w�u �u�u�u�u�N������E  ;�wh{  hY�@ hF�@ �s������ދE�PU�U��U�} ta�E��0��tX�Fuh�  hy�@ h`�@ �5������Ft/�F$;�w&�u �ujS�u�U���R�u�u������� �  +؃E�럋M�IM�M��M��E��0����   �Fuh�  h��@ h��@ ��������FtW�F$;�wN�u �uj S�u��U���R�u�u�X����� �} �?  �u �ujj �u��u��u�u�0����� �  +؃E��p����M�y.}�}�7��uh�  h��@ h��@ �0������E�   �Ft	�F�E�v�Fuh�  h׷@ h��@ ��������E��n ;�v+��   �WU��E�   �@t	�H�M�@�}�v�u �uS�7R�w   ����u �ujSj PR������3ۃ�;}�s��u �uj j �u��u��u�u�=����� �} t(�u �ujj �u��u��u�u������ ��������_^[��]�U����SVW�]�u�CuhH  h��@ h޷@ �������C�@uhI  h>�@ h�@ ��������S�U��[�{ ��uhR  hN�@ hE�@ ��������} u���m��E�E3����E��M�;M�v�}� th[  h}�@ hU�@ �������M���)M;}sh\  h��@ h��@ �m������E��+��} t0�u�uj�uj SV�Z������+3�u�ujWj SV�A������U��E����u�_^[YY]�U��SVW�}�u��Cuh�  h��@ h��@ ��������C��P��Pt���H�{�u���>�} u�S֋ڋ��]+s�+[��{� th�  h�@ h��@ �������C���_^[]�U��U�B�x u3�]�+PP�:����]�U����3�SVW�E��} u3��  �U�B�E��U)U��M�A tu�E�@uh   h�@ h�@ �������U�
�Auh  hA�@ h�@ ��������E��J�Auh  h��@ hH�@ ��������E��J�A �E��U�Bt:�M��@t�U�
�Auh  h�@ h��@ �������E��B$�  �}� )�U�Bu �M�A����u�]�E��(  3��  �]�; u���  �Ct)��@uh[  h�@ h�@ �"�������r�u���3�u��   �E��@��   �U�r�u�M��Aty�M��A tp�Ctj3��E��@uh}  hF�@ h�@ �������Ct�US�U���K�M��E���U��Ct�p�C@t�E�V�E�P�u��a������E��u�E��@t�~�v�Fuh�  hv�@ hM�@ �J������~ ;}�s)}����������E�s��   t�EC�E���S�U���   t)�M��Auh�  h��@ h}�@ ��������M�A�E���   ��   3��E��@uh�  h��@ h��@ �������U���   �J�M�E��U�t�x�֋E��H�E��@u�E��M��At*�M��A t!��   tW�E�P�u��A������E�U�U�}� ��   ��   tM�M�f�y t,�E��x}��uh  hȺ@ hź@ ��������@ �3��U�;�r�   �	�   �3��E��@t�u�u�u��u��u��������-�u�u�u�+���Y3ҊЃ����Q�u�W�u��u���������   t(�M�A t�E3ҊP ���   t�M��@����E��׋փ�����   ��H��Hu�m��M��At8�M�A�E�U�z t�M��AP�U��r�u��������A�u������Y�6�M��At$�E�x t�U��JQ�E��p�u��G������	�u�����Y3҉U��˃��;M�����3�_^[��]Ð�������Ð���QUVWRSPT�q j �q��q�q�q�q�q�q�q�1�_�����LÐ��U��İ�M��u�E�&   �E�   3��M��E��I�{   �{   �E��������]ÐU����SVW�]��}�u��͑����    uh�  h��@ h�@ ������訑����   蝑�����   �C(�E�d�5    ��uh�  h�@ h�@ �������;s(th�  h&�@ h�@ �������E��M��P�A�M�f�f�QS�;����CYt3ɉKRS�SY���A �8u�ujj�P������]��}�u���E�U��R�m ��P�_^[��]Ð��U��Ĭ��@ SVW�����U�E�z�P�UԋMԋ]+Y�]̋E�P�UȋM�9���u3��U�d�    �  �L����M�Aty�=8�@  upj �u�u��������u�>���uA�Eԋ��t8�j�w�3�w�w�<�������t����; u��8�@ �����8�@  �   �U�d�    �  �=8�@  ��   �M�9�����   �uԋ����   �E� �O��3�P�õ@ �Ɗ:
u��t�H:Ju������u�u�E�j�w�3�w�w��������u[���; u��}� tHW����Y�u�Vj j j jh�@ j �E�f�E� P�8�@  ��  Y�U��E�Rh��@ �������$��P����M�Y����  ��E��0�UЃ��M��1�M����E����8  �$���@ ߅@ ��@ Y�@ ��@ ߅@ ߅@ �U�
�����t�'  �Eԋ0���U�W�u��������E��}� u�  ���A �9t
���A �8u+�U�:���r�M�9���v�u�u�ujj�������a�����   ��T�����   �U�W(�M��O,�w0�u��E��0�u�u������S�u�u�������Ef�U�f�P�}�u�u��u�W�u�u�������������   ����A �9u6�}�u0�w�_���Y�؀D t�GR��G@PS����YPSVjj��������{   �{   �{   �Ƌ]ȋM��'�����   �U�:�����   �M�M��E�E��E��U�]�
�K�U�B�Mԋ1���A SUVW�{   �{   �M̻��A �p���_^][��U�:���t{�M�U��B�Mԋ1��}"�U�Bt�Mf�]�f�Y3��U�d�    �^��u�>�M3ۉY���EЉE��؋Eԋ40�����ֵ@ ��th�  h#�@ h��@ �������]Ѕ��u����   �U�d�    _^[��]�U���ܸ �@ �H���f�E� �u�"���Y�E��|�@ �M��E�d�    �E��]�U���ܸL�@ �����E�   �M��} t/f�E� �|�@ �M��M�j �u�׌�����Et	�u�^���Y�E�d�    ��]�    0     w   D T                   <�@  X std::bad_exception  �@                    U���ܸd�@ S�]�P����t�@ �|�@ ����E���U�d�    [��]Ð�   �  ��@ bad_exception * �%�A �%�A �%�A �%�A �%�A �%�A �%�A �% �A �%$�A �%(�A �%,�A �%0�A �%4�A �%8�A �%<�A �%@�A �%D�A �%H�A �%L�A �%P�A �%T�A �%X�A �%\�A �%`�A �%d�A �%h�A �%l�A �%p�A �%t�A �%x�A �%|�A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%��A �%ıA ���%ܱA �%�A �%�A ��                                                                                                                                                                                                                                                                                                                                                                                            Embarcadero RAD Studio 29.0 - Copyright 2022 Embarcadero Technologies, Inc.  @ N@ N@ r@        �Y@                 H�@ L�@ lN@ �O@ �P@ $R@ ��@               Nonshared DATA segment required Cannot run multiple instances of a DLL under WIN32s  i@ @ �@ 7@ �������                                ,�@     ����    <�@     ����@  @         X�@     �����@         P@ �@     p@           |�@     ����       ��@     ��@     �����@         �@ �@ borlndmm hrdir_b.c: LoadLibrary != mmdll borlndmm failed borlndmm @Borlndmm@SysGetMem$qqri @Borlndmm@SysFreeMem$qqrpv @Borlndmm@SysReallocMem$qqrpvi @Borlndmm@SysAllocMem$qqri @Borlndmm@SysRegisterExpectedMemoryLeak$qqrpi @Borlndmm@SysUnregisterExpectedMemoryLeak$qqrpi borlndmm @Borlndmm@HeapAddRef$qqrv @Borlndmm@HeapRelease$qqrv hrdir_b.c: GetMem or FreeMem or ReallocMem from borlndmm failed hrdir_b.c: FATAL!!! memory has been allocated prior to heap redirector hook!                    `@ x@ �@ �@ �@        *)@ �,@ �.@ �1@ l@ p@ T&@ h&@ |&@ �&@ l@ p@ T&@ h&@ |&@ �&@ l@ p@                            �&@                            �&@                             �&@   (                         '@   0                         )'@   8                         L'@   @                         u'@   H                         �'@   P                               X                               `                               h                               p                               x                               �                               �                               �                               �                               �                               �                               �                               �                               �                               �                                                                                                                           0                              @                              `                              �                              �                              �                              �                                                            @                              p                              �                              �                                                             p                              �                                                             �                              �                              `                              �                              p                                                            �                              �                              P	                              0
                              0
                              0
                             Local\FastMM_PID_???????  0123456789ABCDEF The memory manager cannot be changed after it has been used. Cannot Switch Memory Manager   �7@                       	                      
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                2    `  `  `                                                                                                                                                                                               @  �@     allocating handle lock table creating handle lock hlocks handles.c creating global handle lock   ),(((((),(((),#,*((((**##%(*,** &*1*#* * �l�@ t�@ ��@ ��@ ��@ ɣ@ ۣ@ �@  �@ �@ /�@ C�@ R�@ f�@ s�@ �@ ��@ ��@ Ĥ@ Ҥ@ �@ ��@ �@ �@ ,�@ ?�@ c�@ z�@ ��@ ��@ ��@ ĥ@ ӥ@ ߥ@ �@ ��@ �@ $�@ <�@ L�@ f�@ y�@ ��@ ��@ ʦ@ ئ@ �@ ��@ ��@ 
�@ 2   Error 0 Invalid function number No such file or directory Path not found Too many open files Permission denied Bad file number Memory arena trashed Not enough memory Invalid memory block address Invalid environment Invalid format Invalid access code Invalid data Bad address No such device Attempted to remove current directory Not same device No more files Invalid argument Arg list too big Exec format error Cross-device link Too many open files No child processes Inappropriate I/O control operation Executable file in use File too large No space left on device Illegal seek Read-only file system Too many links Broken pipe Math argument Result too large File already exists Possible deadlock Operation not permitted No such process Interrupted function call Input/output error No such device or address Resource temporarily unavailable Block device required Resource busy Not a directory Is a directory  Filename too long Directory not empty Unknown error :  
        creating global stream lock allocating stream lock table creating stream lock strm_locks streams.c              ب@ ٨@ ڨ@ ۨ@ ܨ@ ݨ@ ި@ ߨ@ �@ �@ �@ �@ �@  �@ �@ �@ ��@  �@ �@ �@               �@ �@ #�@ -�@ 6�@ =�@ F�@ M�@ Q�@ U�@ Y�@ ]�@ a�@ e�@ i�@ q�@ z�@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ é@ ǩ@ ˩@ ϩ@ ө@ ש@ ۩@ ߩ@ �@ �@ �@                    ��@ Ч@     �@ �@ �@ ��@        ($v)  .    / : %H:%M:%S %m/%d/%y %A, %B %d, %Y AM PM Monday Tuesday Wednesday Thursday Friday Saturday Sunday Mon Tue Wed Thu Fri Sat Sun January February March April May June July August September October November December Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec C  C     2  �ߡ�Error: system code page access failure; MBCS table not initialized  Assertion failed:  , file  , line   %02d/%02d/%04d %02d:%02d:%02d.%03d          
 
           ����      mJ@            ����   kK@ yK@ Abnormal program termination    LM@ LM@ LM@     No space for copy of command line   No space for copy of command line   DN@ XN@                                                                            �      ��       creating atexit lock                                                                                                                                                                                                                                                                          An exception (%08X) occurred during DllEntryPoint or DllMain in module:
%s    creating thread data lock   Semaphore error                 ����<notype> id->tpName xxtype.cpp tp1 xxtype.cpp tp2 xxtype.cpp tp1->tpName xxtype.cpp tp2->tpName xxtype.cpp IS_STRUC(base->tpMask) xxtype.cpp IS_STRUC(derv->tpMask) xxtype.cpp derv->tpClass.tpcFlags & CF_HAS_BASES xxtype.cpp ((unsigned *)vtablePtr)[-1] == 0 xxtype.cpp <notype> scopeLen >= 0 xxtype.cpp topTypPtr != 0 && IS_STRUC(topTypPtr->tpMask) xxtype.cpp tgtTypPtr != 0 && IS_STRUC(tgtTypPtr->tpMask) xxtype.cpp srcTypPtr == 0 || IS_STRUC(srcTypPtr->tpMask) xxtype.cpp __isSameTypeID(srcTypPtr, tgtTypPtr) == 0 xxtype.cpp tgtTypPtr != 0 && __isSameTypeID(topTypPtr, tgtTypPtr) == 0 xxtype.cpp srcTypPtr xxtype.cpp ((unsigned *)vtablePtr)[-1] == 0 xxtype.cpp addr xxtype.cpp Can't adjust class address (no base class entry found) !"Can't adjust class address (no base class entry found)" xxtype.cpp       ��@     ����8e@         f@ �@                                                                                                                                                                     �   ___CPPdebugHook         �f@                             ����   d�@    Stack Overflow!             �o@                             ����   ��@                      kp@                             ����   ��@                          nv@                             �v@                             ����   \�@      <�@                       ___CPPdebugHook (ctorMask & 0x0100) != 0 || (ctorMask & 0x0020) == 0 xx.cpp (ctorMask & 0x0080) == 0 xx.cpp what? !"what?" xx.cpp what? !"what?" xx.cpp (dtorMask & 0x0080) == 0 xx.cpp what? !"what?" xx.cpp (mfnMask & 0x0080) == 0 xx.cpp what? !"what?" xx.cpp cctrAddr xx.cpp dtorAddr xx.cpp argType xx.cpp __CPPexceptionList xx.cpp xl xx.cpp xdrPtr->xdERRaddr == xl xx.cpp dscPtr->xdERRaddr == errPtr xx.cpp dscPtr->xdHtabAdr == hdtPtr xx.cpp dscPtr->xdArgCopy == 0 xx.cpp (dscPtr->xdMask & TM_IS_PTR) == 0 xx.cpp mask & TM_IS_PTR xx.cpp dscPtr->xdMask & TM_IS_PTR xx.cpp dscPtr->xdTypeID == dscPtr->xdBase xx.cpp hdtPtr->HDcctrAddr xx.cpp dscPtr->xdSize == size xx.cpp xdrPtr && xdrPtr == *xdrLPP xx.cpp bogus context in Local_unwind() !"bogus context in Local_unwind()" xx.cpp std::bad_exception bogus context in _ExceptionHandler() !"bogus context in _ExceptionHandler()" xx.cpp varType->tpClass.tpcFlags & CF_HAS_DTOR xx.cpp varType->tpClass.tpcDtorAddr xx.cpp (vbFlag && (errPtr->ERRcInitDtc >= varType->tpClass.tpcDtorCount)) || (!vbFlag && (errPtr->ERRcInitDtc >= varType->tpClass.tpcNVdtCount)) || flags xx.cpp varType->tpClass.tpcFlags & CF_HAS_DTOR xx.cpp dtorCnt < varCount xx.cpp IS_STRUC(blType->tpMask) xx.cpp IS_STRUC(blType->tpMask) xx.cpp memType xx.cpp memType->tpClass.tpcFlags & CF_HAS_DTOR xx.cpp varType->tpMask & TM_IS_ARRAY xx.cpp varType->tpArr.tpaElemType->tpClass.tpcFlags & CF_HAS_DTOR xx.cpp vdtCount xx.cpp etdCount <= elemCount || elemCount == 0 xx.cpp dtrCount <= vdtCount xx.cpp IS_CLASS(varType->tpMask) xx.cpp ((unsigned *)vftAddr)[-1] == 0 xx.cpp dttPtr->dttFlags & (DTCVF_PTRVAL|DTCVF_RETVAL) xx.cpp dttPtr->dttType->tpMask & TM_IS_PTR xx.cpp dttPtr->dttType->tpPtr.tppBaseType->tpClass.tpcFlags & CF_HAS_DTOR xx.cpp IS_CLASS(dttPtr->dttType->tpMask) && (dttPtr->dttType->tpClass.tpcFlags & CF_HAS_DTOR) xx.cpp dtvtPtr->dttType->tpMask & TM_IS_ARRAY xx.cpp varType->tpClass.tpcFlags & CF_HAS_DTOR xx.cpp elemType->tpClass.tpcFlags & CF_HAS_DTOR xx.cpp varType->tpMask & TM_IS_ARRAY xx.cpp varType->tpMask & TM_IS_PTR xx.cpp bl xx.cpp **BCCxh1 ��@    ����            ����                  غ@     ,�@           �@     ����       �@     ,�@           8�@     ����       <�@         ������@         <�@ �@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             <�         � � ̱         �� ܱ                     � �  � 6� N� \� v� �� �� �� �� Ҳ � �  � � *� 6� H� Z� l� |� �� �� �� �� γ � �� � *� :� J� ^� p� |� �� �� �� ȴ д ܴ � �� � � $� 2� B�     � �  � 6� N� \� v� �� �� �� �� Ҳ � �  � � *� 6� H� Z� l� |� �� �� �� �� γ � �� � *� :� J� ^� p� |� �� �� �� ȴ д ܴ � �� � � $� 2� B�     N� b� p�     N� b� p�     KERNEL32.DLL USER32.DLL   CloseHandle   CreateFileA   CreateFileMappingA    EnterCriticalSection    ExitProcess   FreeEnvironmentStringsW   GetACP    GetCPInfo   GetCurrentProcessId   GetCurrentThreadId    GetEnvironmentStringsW    GetFileType   GetLastError    GetLocalTime    GetModuleFileNameA    GetModuleHandleA    GetOEMCP    GetProcAddress    GetProcessHeap    GetStartupInfoA   GetStdHandle    GetVersion    GetVersionExA   HeapAlloc   HeapFree    InitializeCriticalSection   InterlockedDecrement    InterlockedIncrement    IsDebuggerPresent   LeaveCriticalSection    LoadLibraryA    MapViewOfFile   OpenFileMappingA    RaiseException    RtlUnwind   SetConsoleCtrlHandler   SetFilePointer    SetHandleCount    SetLastError    Sleep   TlsAlloc    TlsFree   TlsGetValue   TlsSetValue   UnmapViewOfFile   VirtualAlloc    VirtualFree   VirtualQuery    WriteFile   EnumThreadWindows   MessageBoxA   wsprintfA                                                                                                                                                 2�          (� ,� 0� �  <�   WinSCP.sv ___CPPdebugHook                                                                                                                                                                                                                                                                                                                                                                                                                                                         �f�Z          (  �
   � �   0 �    �f�Z      �    H �   ` �   x �   � �	   � �
   � �   � �   � �    �     �   8 �   P �   h �   � �   � �   � �   � �   � �   � �   	 �   (	 �   @	 �   X	 �   p	 �   �	 �   �	 �   �	 �    �	 �!   �	 �"    
 �#   
 �$   0
 �%   H
 �&   `
 �'   x
 �(   �
 �,   �
 �-   �
 �.   �
 �/   �
 �0    �1     �2   8 �E   P �F   h �G   � �H   � �I   � �J   � �K   � �L   � �R    �S   ( �T   @ �U   X �V   p �X   � �Y   � �\   � �]   � �^   � �_     �`    �a   0 �b   H �c   ` �d   x �e   � �f   � �g   � �h   � �i   � �j    �k     �l   8 �m   P �n   h �o   � �p   � �q   � �r   � �s   � �t   � �u    �w   ( �x   @ �y   X �z   p �{   � �|   � �}   � �~   � �   � ��     ��    ��   0 ��   H ��   ` ��   x ��   � ��   � ��   � �9  � �:  � �;   �<    �=  8 �>  P �x  h �y  � �z  � �{  � �|  � �}  � �~  � ��   ��  ( ��  @ �  X �  p �  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � ��  � ��   ��  ( ��  @ ��  X ��  p ��  � ��  � ��  � ��  � ��  � ��    ��   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � ��  � �    �    �f�Z    )   �) �( �* �@ � * �X �D* �p �b* �� ��* �� ��* �� ��* �� ��* �� �+ �  �8+ � �f+ �0 ��+ �H ��+ �` ��+ �x ��+ �� �, �� �D, �� �d, �� ��, �� ��, � ��, �  �- �8 �.- �P �^- �h �x- �� ��- �� ��- �� ��- �� �. �� �(. �� �L. � �x. �( ��. �@ ��. �X ��. �p ��. �� �$/ �� �B/ �� �z/ �� ��/ �� �    �f�Z            �    �f�Z               �f�Z         (      �f�Z         8      �f�Z         H      �f�Z         X      �f�Z         h      �f�Z         x      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z               �f�Z               �f�Z         (      �f�Z         8      �f�Z         H      �f�Z         X      �f�Z         h      �f�Z         x      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z               �f�Z               �f�Z         (      �f�Z         8      �f�Z         H      �f�Z         X      �f�Z         h      �f�Z         x      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z               �f�Z               �f�Z         (      �f�Z         8      �f�Z         H      �f�Z         X      �f�Z         h      �f�Z         x      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z         �      �f�Z                �f�Z                �f�Z         (       �f�Z         8       �f�Z         H       �f�Z         X       �f�Z         h       �f�Z         x       �f�Z         �       �f�Z         �       �f�Z         �       �f�Z         �       �f�Z         �       �f�Z         �       �f�Z         �       �f�Z         �       �f�Z         !      �f�Z         !      �f�Z         (!      �f�Z         8!      �f�Z         H!      �f�Z         X!      �f�Z         h!      �f�Z         x!      �f�Z         �!      �f�Z         �!      �f�Z         �!      �f�Z         �!      �f�Z         �!      �f�Z         �!      �f�Z         �!      �f�Z         �!      �f�Z         "      �f�Z         "      �f�Z         ("      �f�Z         8"      �f�Z         H"      �f�Z         X"      �f�Z         h"      �f�Z         x"      �f�Z         �"      �f�Z         �"      �f�Z         �"      �f�Z         �"      �f�Z         �"      �f�Z         �"      �f�Z         �"      �f�Z         �"      �f�Z         #      �f�Z         #      �f�Z         (#      �f�Z         8#      �f�Z         H#      �f�Z         X#      �f�Z         h#      �f�Z         x#      �f�Z         �#      �f�Z         �#      �f�Z         �#      �f�Z         �#      �f�Z         �#      �f�Z         �#      �f�Z         �#      �f�Z         �#      �f�Z         $      �f�Z         $      �f�Z         ($      �f�Z         8$      �f�Z         H$      �f�Z         X$      �f�Z         h$      �f�Z         x$      �f�Z         �$      �f�Z         �$      �f�Z         �$      �f�Z         �$      �f�Z         �$      �f�Z         �$      �f�Z         �$      �f�Z         �$      �f�Z         %      �f�Z         %      �f�Z         (%      �f�Z         8%      �f�Z         H%      �f�Z         X%      �f�Z         h%      �f�Z         x%      �f�Z         �%      �f�Z         �%      �f�Z         �%      �f�Z         �%      �f�Z         �%      �f�Z         �%      �f�Z         �%      �f�Z         �%      �f�Z         &      �f�Z         &      �f�Z         (&      �f�Z         8&      �f�Z         H&      �f�Z         X&      �f�Z         h&      �f�Z         x&      �f�Z         �&      �f�Z         �&      �f�Z         �&      �f�Z         �&      �f�Z         �&      �f�Z         �&      �f�Z         �&      �f�Z         �&      �f�Z         '      �f�Z         '      �f�Z         ('      �f�Z         8'      �f�Z         H'      �f�Z           X'      �f�Z           h'      �f�Z           x'      �f�Z           �'      �f�Z           �'      �f�Z           �'      �f�Z           �'      �f�Z           �'      �f�Z           �'      �f�Z           �'      �f�Z           �'      �f�Z           (      �f�Z           (      �f�Z           ((      �f�Z           8(      �f�Z           H(      �f�Z           X(      �f�Z           h(      �f�Z           x(      �f�Z           �(      �f�Z           �(      �f�Z           �(      �f�Z           �(      �f�Z           �(      �f�Z           �(      �f�Z           �(      �f�Z           �(      �f�Z           )      �f�Z           )      �f�Z           ()      �f�Z           8)      �f�Z           H)      �f�Z           X)      �f�Z           h)      �f�Z           x)      �f�Z           �)      �f�Z           �)      �f�Z           �)      �f�Z           �)      �f�Z           �)      �f�Z           �)      �f�Z       	  �)  �� �          t J          xc R          �g V          $m           Dr v          �v �          �{ ^          � �          � �          ��           �� r          � j          p� &          ��           �� �          8� v          �� �          D� >          �� 4          �� �
          �� 2          �� �          �� P          �� &           � �          � �          �� r          l� �          \� |          �� �          �� �          @ �           � �          d �          H �          � �          �
 �          � �          � R          � �          �& �          @* �           �* �           �+ d          (/ 4          \7 ~          �B :          J           0N &          XU >          �\ �          |c h          �g V          <} �          0� .          `� \          �� p          ,�           @� �          ,� �          Ȳ �          \� �	          �� L          H� �          � 
	           � l          �� �           p� F          ��            �� v           0� *          \� �          �� �          �� �          P� �          �� �          �� �          p� �          H� �           �� �          l� "          �� N          �� X          8 H          � �          t	 �          d �          � �          � �          � �           �           �            � Z          � p          l (          �  l            ! �           �! &           �! �           �" �          `' �           8( (          `, .          �4 p	           > �           F �	          �O �           �P t          V "          ([           ,_ .          \` l          �b R          f �          �g �          �l �           �m p          o >           \o           lp �          0u �          �x �          d} x          ܂ N          ,� D	          p� 4          �� H          � X
          D� �          8� �          ȷ �           �� Z          � �          � r          x�           �� �          \� �          @� �          � D          T� 	          h�           �� �          0� �          0� �          �� :          ,� �          �� �          ��           �� L          �� $          � �           �� �          � D            \          \ �          L �            �          � 2          � :           \          x! Z          �% �          �*           �/           �1 �          P6 :          �: �          l?           |C           �G �          <K �           O �          �Q �           �R �           DS �          �V l          `[ �          X^ �          Ha r          �d            �d A          p l          |�           �� �         l� �          \� �          4� �          �� .          ,� y          �� �          �� �
          �� �          t� c!          � �          � ��         ��	           �
 n�          0�
 �          ��
 �          X�
 0          ��
 s          ��
 �          � ��          4�          L� �          Ԟ �*         �� �          8� ��          �� �         �u �          �� �          t� �          �� �          �* `d          � �	          ̘ �9         ��           �� �         ��           Ȕ n@          8� <           D V C L A L  T A B O U T D I A L O G  T A U T H E N T I C A T E F O R M  T C L E A N U P D I A L O G  T C O N S O L E D I A L O G  T C O P Y D I A L O G  T C O P Y L O C A L D I A L O G  T C O P Y P A R A M C U S T O M D I A L O G  T C O P Y P A R A M P R E S E T D I A L O G  T C O P Y P A R A M S F R A M E  T C R E A T E D I R E C T O R Y D I A L O G  T C U S T O M C O M M A N D D I A L O G  T C U S T O M D I A L O G  T C U S T O M S C P E X P L O R E R F O R M  T E D I T M A S K D I A L O G  T E D I T O R F O R M  T E D I T O R P R E F E R E N C E S D I A L O G  T F I L E F I N D D I A L O G  T F I L E S Y S T E M I N F O D I A L O G  T F U L L S Y N C H R O N I Z E D I A L O G  T G E N E R A T E U R L D I A L O G  T I M P O R T S E S S I O N S D I A L O G  T L I C E N S E D I A L O G  T L O C A T I O N P R O F I L E S D I A L O G  T L O G I N D I A L O G  T M E S S A G E F O R M  T N O N V I S U A L D A T A M O D U L E  T O P E N D I R E C T O R Y D I A L O G  T P R E F E R E N C E S D I A L O G  T P R O G R E S S F O R M  T P R O P E R T I E S D I A L O G  T R E M O T E T R A N S F E R D I A L O G  T R I G H T S F R A M E  T S C P C O M M A N D E R F O R M  T S C P E X P L O R E R F O R M  T S E L E C T M A S K D I A L O G  T S I T E A D V A N C E D D I A L O G  T S Y M L I N K D I A L O G  T S Y N C H R O N I Z E C H E C K L I S T D I A L O G  T S Y N C H R O N I Z E D I A L O G  T S Y N C H R O N I Z E P R O G R E S S F O R M           � H e l p   [   < k o m m a n d o >   [   < k o m m a n d o 2 >   . . .   ] 
     V i s a r   l i s t a   p �   k o m m a n d o n   o m   i n g a   p a r a m e t e r a r   a n g e s . 
     V i s a r   h j � l p   o m   e t t   k o m m a n d o   o m   d e t   a n g e s . 
 a l i a s : 
     m a n 
 e x e m p e l : 
     h e l p 
     h e l p   l s 
 D e x i t 
     S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t . 
 a l i a s : 
     b y e 
 @o p e n   < s i t e > 
 o p e n   s f t p | s c p | f t p [ e s ] | d a v [ s ] | s 3   : / /   [   < u s e r >   [   : p a s s w o r d   ]   @   ]   < h o s t >   [   : < p o r t >   ] 
     E s t a b l i s h e s   c o n n e c t i o n   t o   g i v e n   h o s t .   U s e   e i t h e r   n a m e   o f   t h e   s i t e   o r 
     s p e c i f y   h o s t ,   u s e r n a m e ,   p o r t   a n d   p r o t o c o l   d i r e c t l y . 
 s w i t c h e s : 
     - p r i v a t e k e y = < f i l e >   S S H   p r i v a t e   k e y   f i l e 
     - h o s t k e y = < f i n g e r p r i n t >   F i n g e r p r i n t   o f   s e r v e r   h o s t   k e y   ( S F T P   a n d   S C P   o n l y ) . 
     - c l i e n t c e r t = < f i l e >   T L S / S S L   c l i e n t   c e r t i f i c a t e   f i l e 
     - c e r t i f i c a t e = < f i n g e r p r i n t >   F i n g e r p r i n t   o f   T L S / S S L   c e r t i f i c a t e 
                                           ( F T P S   a n d   W e b D A V S   o n l y ) 
     - p a s s p h r a s e = < p h r >     P r i v a t e   k e y   p a s s p h r a s e 
     - p a s s i v e = o n | o f f         P a s s i v e   m o d e   ( F T P   p r o t o c o l   o n l y ) 
     - i m p l i c i t                     I m p l i c i t   T L S / S S L   ( F T P   p r o t o c o l   o n l y ) 
     - e x p l i c i t                     E x p l i c i t   T L S / S S L   ( F T P   p r o t o c o l   o n l y ) 
     - t i m e o u t = < s e c >           S e r v e r   r e s p o n s e   t i m e o u t 
     - u s e r n a m e = < u s e r >       A n   a l t e r n a t i v e   w a y   t o   p r o v i d e   a   u s e r n a m e 
     - p a s s w o r d = < p a s s w o r d >   A n   a l t e r n a t i v e   w a y   t o   p r o v i d e   a   p a s s w o r d 
     - r a w s e t t i n g s   s e t t i n g 1 = v a l u e 1   s e t t i n g 2 = v a l u e 2   . . . 
                                           C o n f i g u r e s   a n y   s i t e   s e t t i n g s   u s i n g   r a w   f o r m a t 
                                           a s   i n   a n   I N I   f i l e 
     - f i l e z i l l a                   L o a d   < s i t e >   f r o m   F i l e Z i l l a   s i t e   m a n a g e r 
     - n e w p a s s w o r d = < p a s s w o r d >   C h a n g e s   p a s s w o r d   t o   < p a s s w o r d > 
     - p a s s w o r d s f r o m f i l e s   R e a d   a l l   p a s s w o r d s   f r o m   f i l e s 
 e x a m p l e s : 
     o p e n 
     o p e n   s f t p : / / m a r t i n @ e x a m p l e . c o m : 2 2 2 2   - p r i v a t e k e y = m y k e y . p p k 
     o p e n   m a r t i n @ e x a m p l e . c o m 
     o p e n   e x a m p l e . c o m 
 � c l o s e   [   < s e s s i o n >   ] 
     S t � n g e r   s e s s i o n   s p e c i f i c e r a d   m e d   s i t t   n u m m e r .   O m   s e s s i o n s n u m r e t   i n t e   � r 
     s p e c i f i c e r a d ,   s t � n g s   d e n   a k t u e l l a   s e s s i o n e n . 
 e x e m p e l : 
     c l o s e 
     c l o s e   1 
 � s e s s i o n   [   < s e s s i o n >   ] 
     G � r   s e s s i o n e n   s p e c i f i c e r a d   m e d   e t t   n u m m e r   a k t i v .   O m   e t t   s e s s i o n s n u m m e r 
     i n t e   � r   s p e c i f i c e r a d ,   l i s t a s   a n s l u t n a   s e s s i o n e r . 
 e x e m p e l : 
     s e s s i o n 
     s e s s i o n   1 
 ; p w d 
     V i s a r   a k t u e l l   f j � r r k a t a l o g   f � r   d e n   a k t i v a   s e s s i o n e n . 
 � c d   [   < k a t a l o g >   ] 
     � n d r a r   a k t u e l l   k a t a l o g   p �   s e r v e r n   i   d e n   a k t i v a   s e s s i o n e n . 
     O m   e n   k a t a l o g   i n t e   a n g e s ,   a n v � n d s   h e m k a t a l o g e n . 
 e x e m p e l : 
     c d   / h o m e / m a r t i n 
     c d 
 Ul s   [   < d i r e c t o r y >   ] / [   < w i l d c a r d >   ] 
     L i s t s   t h e   c o n t e n t s   o f   s p e c i f i e d   r e m o t e   d i r e c t o r y .   I f   d i r e c t o r y   i s   
     n o t   s p e c i f i e d ,   l i s t s   w o r k i n g   d i r e c t o r y . 
     W h e n   w i l d c a r d   i s   s p e c i f i e d ,   i t   i s   t r e a t e d   a s   s e t   o f   f i l e s   t o   l i s t . 
     O t h e r w i s e ,   a l l   f i l e s   a r e   l i s t e d . 
 a l i a s : 
     d i r 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     l s 
     l s   * . h t m l 
     l s   / h o m e / m a r t i n 
 @ l p w d 
     V i s a r   a k t u e l l   l o k a l   k a t a l o g   ( g � l l e r   f � r   a l l a   s e s s i o n e r ) . 
 J l c d   < k a t a l o g > 
     B y t e r   l o k a l   k a t a l o g   f � r   a l l a   s e s s i o n e r . 
 e x e m p e l : 
     c d   d : \ 
 Bl l s   [   < d i r e c t o r y >   ] \ [   < w i l d c a r d >   ] 
     L i s t s   t h e   c o n t e n t s   o f   s p e c i f i e d   l o c a l   d i r e c t o r y .   I f   d i r e c t o r y   i s   
     n o t   s p e c i f i e d ,   l i s t s   w o r k i n g   d i r e c t o r y . 
     W h e n   w i l d c a r d   i s   s p e c i f i e d ,   i t   i s   t r e a t e d   a s   s e t   o f   f i l e s   t o   l i s t . 
     O t h e r w i s e ,   a l l   f i l e s   a r e   l i s t e d . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     l l s 
     l l s   * . h t m l 
     l l s   d : \ 
 9r m   < f i l e >   [   < f i l e 2 >   . . .   ] 
     R e m o v e s   o n e   o r   m o r e   r e m o t e   f i l e s .   I f   r e m o t e   r e c y c l e   b i n   i s 
     c o n f i g u r e d ,   m o v e s   f i l e   t o   t h e   b i n   i n s t e a d   o f   d e l e t i n g   i t . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     r m   i n d e x . h t m l 
     r m   i n d e x . h t m l   a b o u t . h t m l 
     r m   * . h t m l 
 � r m d i r   < k a t a l o g >   [   < k a t a l o g 2 >   . . .   ] 
     R a d e r a r   e n   e l l e r   f l e r a   f j � r r k a t a l o g e r .   O m   f j � r r p a p p e r s k o r g e n   � r 
   k o n f i g u r e r a d ,   f l y t t a s   k a t a l o g e n   d i t   i s t � l l e t   f � r   a t t   r a d e r a s . 
 e x e m p e l : 
     r m d i r   p u b l i c _ h t m l 
 ?m v   < f i l e >   [   < f i l e 2 >   . . .   ]   [   < d i r e c t o r y > /   ] [   < n e w n a m e >   ] 
     M o v e s   o r   r e n a m e s   o n e   o r   m o r e   r e m o t e   f i l e s .   D e s t i n a t i o n   d i r e c t o r y   o r   n e w 
     n a m e   o r   b o t h   m u s t   b e   s p e c i f i e d .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h   
     s l a s h .   O p e r a t i o n   m a s k   c a n   b e   u s e d   i n s t e a d   o f   n e w   n a m e . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 a l i a s : 
     r e n a m e 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     m v   i n d e x . h t m l   p u b l i c _ h t m l / 
     m v   i n d e x . h t m l   a b o u t . * 
     m v   i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . * 
     m v   p u b l i c _ h t m l / i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . h t m l   / h o m e / m a r t i n / * . b a k 
     m v   * . h t m l   / h o m e / b a c k u p / * . b a k 
 ^c h m o d   < m o d e >   < f i l e >   [   < f i l e 2 >   . . .   ] 
     C h a n g e s   p e r m i s s i o n s   o f   o n e   o r   m o r e   r e m o t e   f i l e s .   M o d e   c a n   b e   s p e c i f i e d 
     a s   t h r e e   o r   f o u r - d i g i t   o c t a l   n u m b e r . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     c h m o d   6 4 4   i n d e x . h t m l   a b o u t . h t m l 
     c h m o d   1 7 0 0   / h o m e / m a r t i n / p u b l i c _ h t m l 
     c h m o d   6 4 4   * . h t m l 
 t l n   < m � l >   < s y m b o l i s k   l � n k > 
     S k a p a r   s y m b o l i s k   f j � r r l � n k . 
 a l i a s : 
     s y m l i n k 
 e x e m p e l : 
     l n   / h o m e / m a r t i n / p u b l i c _ h t m l   w w w 
 D m k d i r   < k a t a l o g > 
     S k a p a r   f j � r r k a t a l o g . 
 e x e m p e l : 
     m k d i r   p u b l i c _ h t m l 
 g e t   < f i l e >   [   [   < f i l e 2 >   . . .   ]   < d i r e c t o r y > \ [   < n e w n a m e >   ]   ] 
     D o w n l o a d s   o n e   o r   m o r e   f i l e s   f r o m   r e m o t e   d i r e c t o r y   t o   l o c a l   d i r e c t o r y . 
     I f   o n l y   o n e   p a r a m e t e r   i s   s p e c i f i e d   d o w n l o a d s   t h e   f i l e   t o   l o c a l   w o r k i n g 
     d i r e c t o r y .   I f   m o r e   p a r a m e t e r s   a r e   s p e c i f i e d ,   a l l   e x c e p t   t h e   l a s t   o n e 
     s p e c i f y   s e t   o f   f i l e s   t o   d o w n l o a d .   T h e   l a s t   p a r a m e t e r   s p e c i f i e s   t a r g e t 
     l o c a l   d i r e c t o r y   a n d   o p t i o n a l l y   o p e r a t i o n   m a s k   t o   s t o r e   f i l e ( s )   u n d e r 
     d i f f e r e n t   n a m e .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h   b a c k s l a s h .   
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
     T o   d o w n l o a d   m o r e   f i l e s   t o   c u r r e n t   w o r k i n g   d i r e c t o r y   u s e   ' . \ '   a s   t h e 
     l a s t   p a r a m e t e r . 
 a l i a s : 
     r e c v ,   m g e t 
 s w i t c h e s : 
     - d e l e t e                     D e l e t e   s o u r c e   r e m o t e   f i l e ( s )   a f t e r   t r a n s f e r 
     - r e s u m e                     R e s u m e   t r a n s f e r   i f   p o s s i b l e   ( S F T P   a n d   F T P   p r o t o c o l s   o n l y ) 
     - a p p e n d                     A p p e n d   f i l e   t o   e n d   o f   t a r g e t   f i l e   ( S F T P   p r o t o c o l   o n l y ) 
     - p r e s e r v e t i m e         P r e s e r v e   t i m e s t a m p 
     - n o p r e s e r v e t i m e     D o   n o t   p r e s e r v e   t i m e s t a m p 
     - s p e e d = < k b p s >         L i m i t   t r a n s f e r   s p e e d   ( i n   K B / s ) 
     - t r a n s f e r = < m o d e >   T r a n s f e r   m o d e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >   S e t s   f i l e   m a s k . 
     - r e s u m e s u p p o r t = < s t a t e >   C o n f i g u r e s   r e s u m e   s u p p o r t . 
                                       P o s s i b l e   v a l u e s   a r e   ' o n ' ,   ' o f f '   o r   t h r e s h o l d 
     - n e w e r o n l y               T r a n s f e r   n e w   a n d   u p d a t e d   f i l e s   o n l y 
     - l a t e s t                     T r a n s f e r   t h e   l a t e s t   f i l e   o n l y 
 e f f e c t i v e   o p t i o n s : 
     c o n f i r m ,   f a i l o n n o m a t c h ,   r e c o n n e c t t i m e 
 e x a m p l e s : 
     g e t   i n d e x . h t m l 
     g e t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . \ 
     g e t   i n d e x . h t m l   a b o u t . h t m l   d : \ w w w \ 
     g e t   p u b l i c _ h t m l / i n d e x . h t m l   d : \ w w w \ a b o u t . * 
     g e t   * . h t m l   * . p n g   d : \ w w w \ * . b a k 
 �p u t   < f i l e >   [   [   < f i l e 2 >   . . .   ]   < d i r e c t o r y > / [   < n e w n a m e >   ]   ] 
     U p l o a d s   o n e   o r   m o r e   f i l e s   f r o m   l o c a l   d i r e c t o r y   t o   r e m o t e   d i r e c t o r y . 
     I f   o n l y   o n e   p a r a m e t e r   i s   s p e c i f i e d   u p l o a d s   t h e   f i l e   t o   r e m o t e   w o r k i n g 
     d i r e c t o r y .   I f   m o r e   p a r a m e t e r s   a r e   s p e c i f i e d ,   a l l   e x c e p t   t h e   l a s t   o n e 
     s p e c i f y   s e t   o f   f i l e s   t o   u p l o a d .   T h e   l a s t   p a r a m e t e r   s p e c i f i e s   t a r g e t 
     r e m o t e   d i r e c t o r y   a n d   o p t i o n a l l y   o p e r a t i o n   m a s k   t o   s t o r e   f i l e ( s )   u n d e r 
     d i f f e r e n t   n a m e .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h   s l a s h .   
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
     T o   u p l o a d   m o r e   f i l e s   t o   c u r r e n t   w o r k i n g   d i r e c t o r y   u s e   ' . / '   a s   t h e 
     l a s t   p a r a m e t e r . 
 a l i a s : 
     s e n d ,   m p u t 
 s w i t c h e s : 
     - d e l e t e                           D e l e t e   s o u r c e   l o c a l   f i l e ( s )   a f t e r   t r a n s f e r 
     - r e s u m e                           R e s u m e   t r a n s f e r   i f   p o s s i b l e   ( S F T P   a n d   F T P   p r o t o c o l s   o n l y ) 
     - a p p e n d                           A p p e n d   f i l e   t o   e n d   o f   t a r g e t   f i l e   ( S F T P   p r o t o c o l   o n l y ) 
     - p r e s e r v e t i m e               P r e s e r v e   t i m e s t a m p 
     - n o p r e s e r v e t i m e           D o   n o t   p r e s e r v e   t i m e s t a m p 
     - p e r m i s s i o n s = < m o d e >   S e t   p e r m i s s i o n s 
     - n o p e r m i s s i o n s             K e e p   d e f a u l t   p e r m i s s i o n s 
     - s p e e d = < k b p s >               L i m i t   t r a n s f e r   s p e e d   ( i n   K B / s ) 
     - t r a n s f e r = < m o d e >         T r a n s f e r   m o d e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >         S e t s   f i l e   m a s k . 
     - r e s u m e s u p p o r t = < s t a t e >   C o n f i g u r e s   r e s u m e   s u p p o r t . 
                                             P o s s i b l e   v a l u e s   a r e   ' o n ' ,   ' o f f '   o r   t h r e s h o l d 
     - n e w e r o n l y                     T r a n s f e r   n e w   a n d   u p d a t e d   f i l e s   o n l y 
     - l a t e s t                           T r a n s f e r   t h e   l a t e s t   f i l e   o n l y 
 e f f e c t i v e   o p t i o n s : 
     c o n f i r m ,   f a i l o n n o m a t c h ,   r e c o n n e c t t i m e 
 e x a m p l e s : 
     p u t   i n d e x . h t m l 
     p u t   - d e l e t e   i n d e x . h t m l   a b o u t . h t m l   . / 
     p u t   - p e r m i s s i o n s = 6 4 4   i n d e x . h t m l   a b o u t . h t m l   / h o m e / m a r t i n / p u b l i c _ h t m l / 
     p u t   d : \ w w w \ i n d e x . h t m l   a b o u t . * 
     p u t   * . h t m l   * . p n g   / h o m e / m a r t i n / b a c k u p / * . b a k 
 �o p t i o n   [   < o p t i o n >   [   < v a l u e >   ]   ] 
     I f   n o   p a r a m e t e r s   a r e   s p e c i f i e d ,   l i s t s   a l l   s c r i p t   o p t i o n s   a n d   t h e i r 
     v a l u e s .   W h e n   o n e   p a r a m e t e r   i s   s p e c i f i e d   o n l y ,   s h o w s   v a l u e   o f   t h e   o p t i o n . 
     W h e n   t w o   p a r a m e t e r s   a r e   s p e c i f i e d   s e t s   v a l u e   o f   t h e   o p t i o n . 
     I n i t i a l   v a l u e s   o f   s o m e   o p t i o n s   a r e   t a k e n   f r o m   a p p l i c a t i o n   c o n f i g u r a t i o n , 
     h o w e v e r   m o d i f i n g   t h e   o p t i o n s   d o e s   n o t   c h a n g e   t h e   a p p l i c a t i o n 
     c o n f i g u r a t i o n . 
 o p t i o n s   a r e : 
     e c h o           o n | o f f 
                       T o g g l e s   e c h o i n g   o f   c o m m a n d   b e i n g   e x e c u t e d . 
                       C o m m a n d s   a f f e c t e d :   a l l 
     b a t c h         o n | o f f | a b o r t | c o n t i n u e 
                       T o g g l e s   b a t c h   m o d e   ( a l l   p r o m p t s   a r e   a u t o m a t i c a l l y   r e p l i e d 
                       n e g a t i v e l y ) .   W h e n   ' o n ' ,   i t   i s   r e c o m m e n d e d   t o   s e t   ' c o n f i r m ' 
                       t o   ' o f f '   t o   a l l o w   o v e r w r i t e s .   W i t h   ' a b o r t ' ,   s c r i p t   i s   a b o r t e d 
                       w h e n   a n y   e r r o r   o c c u r s .   W i t h   ' c o n t i n u e ' ,   a l l   e r r o r s   a r e   i g n o r e d . 
                       R e c o n n e c t   t i m e   i s   a u t o m a t i c a l l y   l i m i t e d   d o   1 2 0 s ,   i f   n o t   l i m i t e d   y e t . 
                       C o m m a n d s   a f f e c t e d :   n e a r l y   a l l 
     c o n f i r m     o n | o f f 
                       T o g g l e s   c o n f i r m a t i o n s   ( o v e r w r i t e ,   e t c . ) . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t 
     r e c o n n e c t t i m e   o f f   |   < s e c > 
                       T i m e   l i m i t   i n   s e c o n d s   t o   t r y   r e c o n n e c t i n g   b r o k e n   s e s s i o n s . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   s y n c h r o n i z e ,   k e e p u p t o d a t e 
     f a i l o n n o m a t c h   o n | o f f 
                       W h e n   ' o n ' ,   c o m m a n d s   f a i l   w h e n   f i l e   m a s k   m a t c h e s   n o   f i l e s . 
                       W h e n   ' o f f ' ,   c o m m a n d s   d o   n o t h i n g   w h e n   f i l e   m a s k   m a t c h e s   n o   f i l e s . 
                       C o m m a n d s   a f f e c t e d :   g e t ,   p u t ,   r m ,   m v ,   c h m o d ,   l s ,   l l s 
 e x a m p l e s : 
     o p t i o n 
     o p t i o n   b a t c h 
     o p t i o n   c o n f i r m   o f f 
 As y n c h r o n i z e   l o c a l | r e m o t e | b o t h   [   < l o k a l   k a t a l o g >   [   < f j � r r k a t a l o g >   ]   ] 
     N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' l o c a l '   s y n k r o n i s e r a s   l o k a l   k a t a l o g   m e d 
     f j � r r k a t a l o g .   N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' r e m o t e '   s y n k r o n i s e r a s   f j � r r k a t a l o g 
     m e d   l o k a l   k a t a l o g .   N � r   d e n   f � r s t a   p a r a m e t e r n   � r   ' b o t h '   s y n k r o n i s e r a s 
     k a t a l o g e r n a   m o t   v a r a n d r a . 
     N � r   k a t a l o g e r   i n t e   s p e c i f i c e r a s ,   s y n k r o n i s e r a s   a k t u e l l 
     k a t a l o g . 
     O B S :   � v e r s k r i v n i n g s b e k r � f t e l s e r   � r   a l l t i d   a v   f � r   k o m m a n d o t . 
 v � x l a r : 
     - p r e v i e w                           F � r h a n d s g r a n s k a   � n d r i n g a r ,   s y n k r o n i s e r a r   i n t e 
     - d e l e t e                             T a   b o r t   f � r � l d r a d e   f i l e r 
     - m i r r o r                             S p e g e l l � g e   ( s y n k r o n i s e r a r   f � r � l d r a d e   f i l e r   o c k s � ) . 
                                               I g n o r e r a s   m e d   ' b o t h ' . 
     - c r i t e r i a = < k r i t e r i e r >   J � m f � r e l s e k r i t e r i e r .   M � j l i g a   v � r d e n   � r   ' n o n e ' ,   ' t i m e ' , 
                                               ' s i z e '   o c h   ' e i t h e r ' .   I g n o r e r a s   m e d   ' b o t h ' - l � g e . 
     - p e r m i s s i o n s = < l � g e >     A n g e   r � t t i g h e t e r 
     - n o p e r m i s s i o n s               B e h � l l   s t a n d a r d r � t t i g h e t e r 
     - s p e e d = < k b p s >               B e g r � n s a   � v e r f � r i n g s h a s t i g h e t 
     - t r a n s f e r = < l � g e >           � v e r f � r i n g s l � g e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >           A n g e   f i l m a s k . 
     - r e s u m e s u p p o r t = < t i l l s t � n d >   K o n f i g u r e r a r   � t e r u p p t a g n i n g s s t � d . 
                                               M � j l i g a   v � r d e n   � r   ' o n ' ,   ' o f f '   e l l e r   t r � s k e l 
 e f f e k t i v a   a l t e r n a t i v : 
     r e c o n n e c t t i m e 
 e x e m p e l : 
     s y n c h r o n i z e   r e m o t e   - d e l e t e 
     s y n c h r o n i z e   b o t h   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 Sk e e p u p t o d a t e   [   < l o c a l   d i r e c t o r y >   [   < r e m o t e   d i r e c t o r y >   ]   ] 
     W a t c h e s   f o r   c h a n g e s   i n   l o c a l   d i r e c t o r y   a n d   r e f l e c t s   t h e m   o n   r e m o t e   o n e . 
     W h e n   d i r e c t o r i e s   a r e   n o t   s p e c i f i e d ,   c u r r e n t   w o r k i n g   d i r e c t o r i e s   a r e 
     s y n c h r o n i z e d .   T o   s t o p   w a t c h i n g   f o r   c h a n g e s   p r e s s   C t r l - C . 
     N o t e :   O v e r w r i t e   c o n f i r m a t i o n s   a r e   a l w a y s   o f f   f o r   t h e   c o m m a n d . 
 s w i t c h e s : 
     - d e l e t e                           D e l e t e   o b s o l e t e   f i l e s 
     - p e r m i s s i o n s = < m o d e >   S e t   p e r m i s s i o n s 
     - n o p e r m i s s i o n s             K e e p   d e f a u l t   p e r m i s s i o n s 
     - s p e e d = < k b p s >               L i m i t   t r a n s f e r   s p e e d   ( i n   K B / s ) 
     - t r a n s f e r = < m o d e >         T r a n s f e r   m o d e :   b i n a r y ,   a s c i i ,   a u t o m a t i c 
     - f i l e m a s k = < m a s k >         S e t s   f i l e   m a s k . 
     - r e s u m e s u p p o r t = < s t a t e >   C o n f i g u r e s   r e s u m e   s u p p o r t . 
                                             P o s s i b l e   v a l u e s   a r e   ' o n ' ,   ' o f f '   o r   t h r e s h o l d 
 e f f e c t i v e   o p t i o n s : 
     r e c o n n e c t t i m e 
 e x a m p l e s : 
     k e e p u p t o d a t e   - d e l e t e 
     k e e p u p t o d a t e   d : \ w w w   / h o m e / m a r t i n / p u b l i c _ h t m l 
 Wc a l l   < K o m m a n d o > 
     M e d   S F T P   o c h   S C P   p r o t o k o l l e n ,   k � r s   g o d t y c k l i g t   f j � r r s k a l s k o m m a n d o . 
     O m   a k t u e l l   s e s s i o n   i n t e   t i l l � t e r   k � r n i n g   a v   g o d t y c k l i g   f j � r r k o m m a n d o 
     s k i l d a   s k a l s e s s i o n e r   k o m m e r   a t t   � p p n a s   a u t o m a t i s k t . 
     O m   F T P   p r o t o k o l l ,   k � r   e t t   p r o t o k o l l k o m m a n d o . 
     K o m m a n d o t   k a n   i n t e   k r � v a   a n v � n d a r i n p u t . 
 a l i a s : 
     ! 
 e x e m p e l : 
     c a l l   t o u c h   i n d e x . h t m l 
 ] e c h o   < m e d d e l a n d e > 
     S k r i v e r   m e d d e l a n d e   t i l l   s k r i p t u t d a t a . 
 e x e m p e l : 
     e c h o   S t a r t i n g   u p l o a d . . . 
 Y s t a t   < f i l > 
     H � m t a r   o c h   l i s t a r   a t t r i b u t   f � r   a n g i v e n   f j � r r f i l . 
 e x e m p e l : 
     s t a t   i n d e x . h t m l 
 a c h e c k s u m   < a l g >   < f i l e > 
     C a l c u l a t e s   c h e c k s u m   o f   r e m o t e   f i l e . 
 e x a m p l e : 
     c h e c k s u m   s h a - 1   i n d e x . h t m l 
 (c p   < f i l e >   [   < f i l e 2 >   . . .   ]   [   < d i r e c t o r y > /   ] [   < n e w n a m e >   ] 
     D u p l i c a t e s   o n e   o r   m o r e   r e m o t e   f i l e s .   D e s t i n a t i o n   d i r e c t o r y   o r   n e w 
     n a m e   o r   b o t h   m u s t   b e   s p e c i f i e d .   D e s t i n a t i o n   d i r e c t o r y   m u s t   e n d   w i t h 
     s l a s h .   O p e r a t i o n   m a s k   c a n   b e   u s e d   i n s t e a d   o f   n e w   n a m e . 
     F i l e n a m e   c a n   b e   r e p l a c e d   w i t h   w i l d c a r d   t o   s e l e c t   m u l t i p l e   f i l e s . 
 e f f e c t i v e   o p t i o n : 
     f a i l o n n o m a t c h 
 e x a m p l e s : 
     c p   i n d e x . h t m l   p u b l i c _ h t m l / 
     c p   i n d e x . h t m l   a b o u t . * 
     c p   i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . * 
     c p   p u b l i c _ h t m l / i n d e x . h t m l   p u b l i c _ h t m l / a b o u t . h t m l   / h o m e / m a r t i n / * . b a k 
     c p   * . h t m l   / h o m e / b a c k u p / * . b a k 
             
 C O R E _ E R R O R " V � r d n y c k e l n   k u n d e   i n t e   v e r i f i e r a s !  A n s l u t n i n g   m i s s l y c k a d e s .  A v s l u t a d   a v   a n v � n d a r e n .  T a p p a d   a n s l u t n i n g . # K a n   i n t e   h i t t a   k o m m a n d o t s   r e t u r k o d . G K o m m a n d o t   ' % s ' 
 m i s s l y c k a d e s   m e d   r e t u r k o d   % d   o c h   f � l j a n d e   f e l m e d d e l a n d e . ) K o m m a n d o t   m i s s l y c k a d e s   m e d   r e t u r k o d e n   % d . 7 K o m m a n d o t   ' % s '   m i s s l y c k a d e s   m e d   o g i l t i g   u t m a t n i n g   ' % s ' . = F e l   u p p s t o d   n � r   n a m n e t   p �   a k t u e l l   f j � r r k a t a l o g   s k u l l e   h � m t a s . | F e l   u p p s t o d   n � r   s t a r t m e d d e l a n d e   h o p p a d e s   � v e r .   D i t t   s k a l   � r   a n t a g l i g e n   i n k o m p a t i b e l t   m e d   a p p l i k a t i o n e n   ( B A S H   r e k o m m e n d e r a s ) . ) F e l   u p p s t o d   n � r   k a t a l o g   b y t t e s   t i l l   ' % s ' .     ) F e l   u p p s t o d   n � r   l i s t n i n g   a v   k a t a l o g   ' % s ' . % O v � n t a d   k a t a l o g l i s t n i n g   v i d   r a d   ' % s ' . # F e l a k t i g   r � t t i g h e t s b e s k r i v n i n g   ' % s ' ; F e l   u p p s t o d   n � r   d e n   a l l m � n n a   k o n f i g u r a t i o n e n   s k u l l e   r e n s a s .   F e l   v i d   r e n s n i n g   a v   c a c h e m i n n e t . 1 F e l   u p p s t o d   n � r   f i l e n   m e d   s l u m p t a l s f r � n   r e n s a d e s . - F e l   u p p s t o d   n � r   c a c h a d e   v � r d n y c k l a r   r e n s a d e s . Q F e l   u p p s t o d   n � r   v a r i a b e l   i n n e h � l l a n d e   r e t u r k o d   a v   s e n a s t e   k o m m a n d o   s k u l l e   h i t t a s . 0 F e l   u p p s t o d   n � r   a n v � n d a r g r u p p e r   s k u l l e   s l � s   u p p . " F i l   e l l e r   k a t a l o g   ' % s '   f i n n s   i n t e . ) K a n   i n t e   h i t t a   a t t r i b u t e n   f � r   f i l e n   ' % s ' .  K a n   i n t e   � p p n a   f i l e n   ' % s ' . ( F e l   u p p s t o d   n � r   f i l e n   ' % s '   s k u l l e   l � s a s . 3 A l l v a r l i g t   f e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l e n   ' % s ' . 0 F i l k o p i e r i n g e n   t i l l   f j � r r k a t a l o g e n   m i s s l y c k a d e s .   0 F i l k o p i e r i n g e n   f r � n   f j � r r k a t a l o g e n   m i s s l y c k a d e s . % S C P   p r o t o k o l l f e l :   O v � n t a d   r a d b r y t n i n g & S C P   p r o t o k o l l f e l :   F e l a k t i g t   t i d s f o r m a t 2 S C P   p r o t o k o l l f e l :   F e l a k t i g   c o n t r o l   r e c o r d   ( % s ;   % s ) # K o p i e r i n g   a v   f i l   ' % s '   m i s s l y c k a d e s . 1 S C P   p r o t o k o l l f e l :   F e l a k t i g t   f i l b e s k r i v n i n g s f o r m a t  ' % s '   � r   i n g e n   k a t a l o g ! ( F e l   u p p s t o d   n � r   k a t a l o g e n   ' % s '   s k a p a d e s .  K a n   i n t e   s k a p a   f i l e n   ' % s ' . * F e l   u p p s t o d   v i d   s k r i v n i n g   t i l l   f i l e n   ' % s ' . * K a n   i n t e   s � t t a   a t t r i b u t e n   t i l l   f i l e n   ' % s ' . + F e l m e d d e l a n d e   m o t t a g e t   f r � n   f j � r r s i d a :   ' % s ' " F e l   v i d   b o r t t a g n i n g   a v   f i l e n   ' % s ' . 7 F e l   u p p s t o d   v i d   l o g g n i n g   o c h   d e n   h a r   d � r f � r   s t � n g t s   a v .  K a n   i n t e   � p p n a   l o g g f i l e n   ' % s ' . 0 F e l   u p p s t o d   n � r   f i l e n   ' % s '   b y t t e   n a m n   t i l l   ' % s ' .     F i l e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . $ K a t a l o g e n   m e d   n a m n   ' % s '   f i n n s   r e d a n . 2 F e l   u p p s t o d   v i d   b y t e   a v   k a t a l o g   t i l l   h e m k a t a l o g e n . ' F e l   u p p s t o d   v i d   r e n s n i n g   a v   a l l a   a l i a s .   ; F e l   u p p s t o d   n � r   n a t i o n e l l a   a n v � n d a r v a r i a b l e r   s k u l l e   r e n s a s . ! O v � n t a d   i n d a t a   f r � n   s e r v e r n :   ' % s ' ( F e l   u p p s t o d   n � r   I N I - f i l e n   s k u l l e   r e n s a s .   6 A u t e n t i s e r i n g s l o g g   ( s e   s e s s i o n s l o g g   f � r   d e t a l j e r ) : 
 % s 
  A u t e n t i s e r i n g   m i s s l y c k a d e s . # A n s l u t n i n g e n   h a r   o v � n t a t   a v s l u t a t s . 1 F e l   u p p s t o d   n � r   n y c k e l n   s p a r a d e s   t i l l   f i l e n   ' % s ' .   ) S e r v e r n   s k i c k a d e   k o m m a n d o t   s l u t s t a t u s   % d . < S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g   m e d d e l a n d e t y p   v i d   s v a r   ( % d ) .   I S F T P - s e r v e r n s   v e r s i o n   ( % d )   s t � d s   i n t e .   V e r s i o n e r   s o m   s t � d s   � r   % d   t i l l   % d . E S F T P   p r o t o k o l l v a r n i n g :   F e l a k t i g t   m e d d e l a n d e n u m m e r   % d   ( f � r v � n t a d e   % d ) .  O v � n t a d   O K   r e s p o n s .  O v � n t a d   E O F   r e s p o n s . ! F i l e n   e l l e r   k a t a l o g e n   f i n n s   i n t e .  � t k o m s t   n e k a d . . A l l m � n t   f e l   ( s e r v e r n   b o r d e   g e   f e l b e s k r i v n i n g ) . J D � l i g t   m e d d e l a n d e   ( D � l i g t   f o r m a t e r a t   p a k e t   e l l e r   i n k o m p a t i b e l t   p r o t o k o l l ) .  I n g e n   a n s l u t n i n g .  F � r l o r a d   a n s l u t n i n g .   S e r v e r n   s t � d e r   i n t e   o p e r a t i o n e n . - % s 
 F e l k o d :   % d 
 F e l m e d d e l a n d e   f r � n   s e r v e r % s :   % s  O k � n d   s t a t u s k o d . ' F e l   v i d   l � s n i n g   a v   s y m b o l i s k   l � n k   ' % s ' . 4 S e r v e r n   r e t u r n e r a d e   t o m   l i s t n i n g   f � r   k a t a l o g e n   ' % s ' . 6 M o t t o g   S S H _ F X P _ N A M E   p a k e t   m e d   n o l l   e l l e r   f l e r a   p o s t e r .   + K a n   i n t e   f �   d e n   v e r k l i g a   s � k v � g e n   f � r   ' % s ' . ) K a n   i n t e   � n d r a   e g e n s k a p e r   f � r   f i l e n   ' % s ' . F K a n   i n t e   i n i t i a l i s e r a   S F T P - p r o t o k o l l e t .   K � r   v � r d d a t o r n   e n   S F T P - s e r v e r ? " K a n   i n t e   l � s a   t i d s z o n s i n f o r m a t i o n .  K a n   i n t e   s k a p a   f j � r r f i l   ' % s ' .  K a n   i n t e   � p p n a   f j � r r f i l   ' % s ' .  K a n   i n t e   s t � n g a   f j � r r f i l   ' % s ' .  ' % s '   � r   i n t e   e n   f i l ! � � v e r f � r i n g e n   l y c k a d e s   s l u t f � r a ,   m e n   t e m p o r � r   � v e r f � r i n g s f i l   ' % s '   k u n d e   i n t e   b y t a   n a m n   t i l l   m � l f i l   ' % s ' .   O m   p r o b l e m e t   k v a r s t � r ,   p r o v a   m e d   a t t   s l �   a v   f i l � v e r f � r i n g e n s   � t e r u p p t a - f u n k t i o n  K a n   i n t e   s k a p a   l � n k   ' % s ' .  O g i l t i g t   k o m m a n d o   ' % s ' .  I n g e n 4 ' % s '   � r   i n g e n   t i l l � t e n   f i l r � t t i g h e t   i   o k t a l t   f o r m a t . 5 S e r v e r n   k r � v e r   e t t   e j   s t � t t   s l u t - p � - r a d   s e k v e n s   ( % s ) .  O k � n d   f i l t y p   ( % d )  O g i l t i g t   v e r k t y g .   % S � k v � g e n   f i n n s   i n t e   e l l e r   � r   o g i l t i g .  F i l e n   f i n n s   r e d a n . R F i l e n   l i g g e r   p �   e n   e n h e t   s o m   e n d a s t   s t � d e r   l � s n i n g ,   e l l e r   e n h e t e n   � r   s k r i v s k y d d a d .   D e t   f i n n s   i n g e t   m e d i a   i   e n h e t e n . * F e l   u p p s t o d   v i d   a v k o d n i n g   a v   U T F - 8   s t r � n g . < F e l   u p p s t o d   v i d   k � r n i n g   a v   e g e t   k o m m a n d o   ' % s '   p �   f i l e n   ' % s ' .  K a n   i n t e   l a d d a   l o c a l e   % d . + M o t t o g   e j   k o m p l e t t a   d a t a p a k e t   f � r e   f i l s l u t . 8 F e l   u p p s t o d   v i d   b e r � k n i n g   a v   s t o r l e k   f � r   k a t a l o g e n   ' % s ' . L M o t t o g   e t t   f � r   s t o r t   ( % d   B )   S F T P   p a k e t .   M a x i m a l t   s t � d d   p a k e t s t o r l e k   � r   % d   B . � K a n   i n t e   k � r a   S C P   f � r   a t t   s t a r t a   � v e r f � r i n g .   K o n t r o l l e r a   a t t   S C P   � r   i n s t a l l e r a t   p �   s e r v e r n   o c h   a t t   s � k v � g e n   � r   i n k l u d e r a d   i   P A T H .   D u   k a n   o c k s �   p r o v a   S F T P   i s t � l l e t   f � r   S C P .  P l a t s p r o f i l e n   ' % s '   f i n n s   r e d a n . , F e l   u p p s t o d   v i d   f l y t t   a v   f i l   ' % s '   t i l l   ' % s ' . x % s 
   
 F e l e t   o r s a k a s   n o r m a l t   a v   e t t   m e d d e l a n d e   f r � n   e t t   i n l o g g n i n g s s k r i p t   ( s o m   . p r o f i l e ) .   M e d d e l a n d e t   k a n   s t a r t a   m e d   " % s " . � * * � v e r f � r i n g   a v   f i l   ' % s '   l y c k a d e s ,   m e n   f e l   u p p s t o d   v i d   i n s t � l l n i n g   a v   r � t t i g h e t e r   o c h / e l l e r   t i d s s t � m p e l . * * 
 
 O m   p r o b l e m e t   k v a r s t � r ,   s t � n g   a v   a n g e   r � t t i g h e t e r   e l l e r   b e v a r a   t i d s s t � m p e l .   A l t e r n a t i v e t   k a n   d u   a k t i v e r a   a l t e r n a t i v e t   ' I g n o r e r a   r � t t i g h e t s f e l ' .  O g i l t i g   � t k o m s t   t i l l   m i n n e t .   2 D e t   f i n n s   i n g e n   l e d i g t   u t r y m m e   k v a r   i   f i l s y s t e m e t . t O p e r a t i o n e n   k a n   i n t e   s l u t f � r a s   p �   g r u n d   a v   a t t   d e t   s k u l l e   m e d f � r a   a t t   a n v � n d a r e n s   l a g r i n g s - q u o t a   s k u l l e   � v e r s k r i d a s . $ P r i n c i p a l   ( % s )   � r   o k � n t   f � r   s e r v e r n . 0 F e l   u p p s t o d   v i d   k o p i e r i n g   a v   f i l   ' % s '   t i l l   ' % s ' . ( O a v s l u t a t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . $ O k � n t   m � n s t e r   ' % s '   v i d   b � r j a n   a v   % d . V K a n   i n t e   k o m b i n e r a   f i l n a m n s m � n s t e r   ( b � r j a r   v i d   % d )   m e d   f i l l i s t m � n s t e r   ( b � r j a r   v i d   % d ) .  O k � n t   k o m m a n d o   ' % s ' . 0 T v e t y d i g t   k o m m a n d o   ' % s ' .   M � j l i g   m a t c h n i n g   � r :   % s $ P a r a m e t e r   s a k n a s   f � r   k o m m a n d o t   ' % s ' . ( F � r   m � n g a   p a r a m e t r a r   f � r   k o m m a n d o t   ' % s ' .          I n g e n   s e s s i o n .  O g i l t i g t   s e s s i o n s n u m m e r   ' % s ' .  O k � n t   a l t e r n a t i v   ' % s ' . % O k � n t   v � r d e   ' % s '   f � r   a l t e r n a t i v   ' % s ' . ( K a n   i n t e   b e s t � m m a   s t a t u s   p �   s o c k e t   ( % d ) . � F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' .   E f t e r   � t e r u p p t a g e n   f i l � v e r f � r i n g   m � s t e   b e f i n t l i g   m � l f i l   t a s   b o r t .   O m   d u   i n t e   h a   r � t t i g h e t e r   a t t   t a   b o r t   m � l f i l ,   m � s t e   d u   a v a k t i v e r a   � t e r u p p t a g n i n g   a v   f i l � v e r f � r i n g . 5 F e l   u p p s t o d   v i d   a v k o d n i n g   a v   S F T P   p a k e t   ( % d ,   % d ,   % d ) . 1 O g i l t i g t   n a m n   ' % s ' .   N a m n   k a n   i n t e   i n n e h � l l a   ' % s ' . @ F i l e n   k u n d e   i n t e   � p p n a s   f � r   a t t   d e n   � r   l � s t   a v   e n   a n n a n   p r o c e s s .  K a t a l o g e n   � r   i n t e   t o m . + D e n   s p e c i f i c e r a d e   f i l e n   � r   i n t e   e n   k a t a l o g .  F i l n a m n e t   � r   i n t e   g i l t i g t . ( F � r   m � n g a   s y m b o l i s k a   l � n k a r   a n t r � f f a d e s .  F i l e n   k a n   i n t e   t a s   b o r t . p E n   a v   p a r a m e t r a r n a   v a r   u t a n f � r   i n t e r v a l l e t ,   e l l e r   p a r a m e t r a r n a   s o m   s p e c i f i c e r a d e s   k a n   i n t e   a n v � n d a s   t i l l s a m m a n s . V D e n   s p e c i f i c e r a d e   f i l e n   v a r   e n   k a t a l o g ,   i   e n   k o n t e x t   d � r   e n   k a t a l o g   i n t e   k a n   a n v � n d a s .  L � s   f � r   b y t e i n t e r v a l l   k r o c k a d e .    L � s   f � r   b y t e i n t e r v a l l   n e k a d e s . P E n   o p e r a t i o n   f � r s � k t e   g � r a s   p �   e n   f i l   s o m   h a r   e n   v � n t a n d e   b o r t t a g n i n g s o p e r a t i o n . F F i l e n   � r   k o r r u p t ;   e n   k o n t r o l l   a v   i n t e g r i t e t e n   i   f i l s y s t e m e t   b � r   k � r a s . ? F i l   ' % s '   i n n e h � l l e r   i n t e   d e n   p r i v a t a   n y c k e l n   i   e t t   k � n t   f o r m a t . e * * D e n   p r i v a t a   n y c k e l f i l e n   ' % s '   i n n e h � l l e r   n y c k e l n   i   f o r m a t e t   % s .   W i n S C P   s t � d e r   e n d a s t   P u T T Y - f o r m a t . * * H D e n   p r i v a t a   n y c k e l f i l e n   ' % s '   i n n e h � l l e r   n y c k e l   i   f � r � l d r a t   S S H - 1 - f o r m a t . � K a n   i n t e   s k r i v a   � v e r   f j � r r f i l e n   ' % s ' . $ $ 
 
 T r y c k   ' T a   b o r t '   f � r   a t t   t a   b o r t   f i l e n   o c h   s k a p a   e n   n y   i   s t � l l e t   f � r   a t t   s k r i v a   � v e r   d e n . $ $  & T a   b o r t = F e l   u p p s t o d   v i d   k o n t r o l l   a v   l e d i g t   u t r y m m e   f � r   s � k v � g e n   ' % s ' . S K a n   i n t e   h i t t a   l e d i g   l o k a l   l i s t n i n g s p o r t n u m m e r   f � r   t u n n e l   i   i n t e r v a l l e t   % d   t i l l   % d . * K a n   i n t e   u t f � r a   n � t v e r k s h � n d e l s e   ( f e l   % d ) . / S e r v e r n   a v s l u t a d e   o v � n t a t   n � t v e r k s a n s l u t n i n g e n . 1 F e l   u p p s t o d   n � r   a n s l u t n i n g e n   s k u l l e   t u n n l a s . 
   
 % s 9 F e l   u p p s t o d   n � r   k o n t r o l l s u m m a n   b e r � k n a d e s   f � r   f i l e n   ' % s ' .  I n t e r n t   f e l   % s   ( % s ) .  O p e r a t i o n e n   s t � d s   i n t e .    � t k o m s t   n e k a d . ' F r � g a r   e f t e r   a u t e n t i s e r i n g s u p p g i f t e r . . . $ O g i l t i g t   s v a r   t i l l   % s   k o m m a n d o   ' % s ' .    O k � n d   v � x e l   ' % s ' . ) F e l   u p p s t o d   v i d   � v e r f � r i n g   a v   f i l e n   ' % s ' .  K a n   i n t e   k � r a   ' % s ' .  F i l e n   ' % s '   h i t t a d e s   i n t e . . E t t   f e l   u p p s t o d   n � r   d o k u m e n t e t   s k u l l e   s t � n g a s . % ' % s '   � r   i n g e n   g i l t i g   h a s t i g h e t s g r � n s .  C e r t i f i k a t k e d j a n   � r   f � r   l � n g .  C e r t i f i k a t   h a r   u p p h � r t .   C e r t i f i k a t   � r   � n n u   i n t e   g i l t i g t .  C e r t i f i k a t   a v v i s a t .  C e r t i f i k a t   s i g n a t u r f e l .  C e r t i f i k a t   e j   s � k e r t .    S j � l v s i g n e r a t   c e r t i f i k a t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - t i l l   f � l t . , F o r m a t   f e l   i   c e r t i f i k a t e t s   g i l t i g - f r � n   f � l t .  O g i l t i g   C A   c e r t i f i k a t .  E j   s t � t t   c e r t i f i k a t   � n d a m � l . 5 N y c k e l a n v � n d n i n g   i n k l u d e r a r   i n t e   c e r t i f i k a t s i g n e r i n g . , B e g r � n s n i n g a r   f � r   s � k v � g s l � n g d e n   � v e r s k r i d s . + S j � l v s i g n e r a t   c e r t i f i k a t   i   c e r t i f i k a t k e d j a . 6 D e t   g � r   i n t e   a t t   a v k o d a   u t f � r d a r e n s   o f f e n t l i g a   n y c k e l . 3 D e t   g � r   i n t e   a t t   d e k r y p t e r a   c e r t i f i k a t e t s   s i g n a t u r . + D e t   g � r   i n t e   a t t   f �   u t f � r d a r e n s   c e r t i f i k a t . 2 D e t   g � r   i n t e   a t t   h � m t a   l o k a l t   u t f � r d a t   c e r t i f i k a t . 3 D e t   g � r   i n t e   a t t   v e r i f i e r a   d e t   f � r s t a   c e r t i f i k a t e t . % O k � n t   f e l   v i d   k o n t r o l l   a v   c e r t i f i k a t . 6 F e l e t   i n t r � f f a d e   p �   e t t   d j u p   a v   % d   i   c e r t i f i k a t k e d j a n .      M a s k e n   � r   o g i l t i g   n � r a   ' % s ' . � S e r v e r n   k a n   i n t e   � p p n a   a n s l u t n i n g   i   a k t i v t   l � g e .   O m   d u   s i t t e r   b a k o m   e n   N A T - r o u t e r ,   k a n   d u   b e h � v a   a n g e   e n   e x t e r n   I P - a d r e s s .   A l t e r n a t i v t ,   � v e r v � g a   a t t   b y t a   t i l l   p a s s i v t   l � g e . ( F e l   u p p s t o d   v i d   b o r t t a g n i n g   a v   f i l   ' % s ' . ? O g i l t i g t   v � r d e   p �   v � x e l   ' % s ' .   G i l t i g a   v � r d e n   � r   ' o n '   o c h   ' o f f ' .   0 K a n   i n t e   � p p n a   w e b b p l a t s k a t a l o g   e l l e r   a r b e t s y t a . ) N � t v e r k s f e l :   I n g e   v � g   t i l l   v � r d   " % H O S T % " . 2 N � t v e r k s f e l :   M j u k v a r a   o r s a k a d e   a v b r u t e n   a n s l u t n i n g  V � r d   " % H O S T % "   f i n n s   i n t e . 0 I n k o m m a n d e   p a k e t   v a r   f � r v a n s k a t   v i d   d e k r y p t e r i n g U % s 
 
 H j � l p   o s s   a t t   f � r b � t t r a   W i n S C P   g e n o m   a t t   r a p p o r t e r a   f e l   p �   W i n S C P : s   s u p p o r t f o r u m . - F e l   v i d   a v k o d n i n g   a v   T L S / S S L - c e r t i f i k a t   ( % s ) .  C O R E _ C O N F I R M A T I O N M V � r d e n   k o m m u n i c e r a r   i n t e   u n d e r   % d   s e k u n d e r . 
 
 V � n t a   y t t e r l i g a r e   % 0 : d   s e k u n d e r ?    & L � s e n o r d   f � r   n y c k e l n   ' % s ' : # F i l e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ' K a t a l o g e n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ?    c h i f f e r  k l i e n t - t i l l - s e r v e r   c h i f f e r  s e r v e r - t i l l - k l i e n t   c h i f f e r � * * V i l l   d u   � t e r u p p t a   f i l � v e r f � r i n g e n ? * * 
 
 M � l k a t a l o g e n   i n n e h � l l e r   d e l v i s   � v e r f � r d   f i l   ' % s ' . 
 
 O B S : S v a r a   ' N e j '   t a r   b o r t   d e l v i s   � v e r f � r d   f i l   o c h   s t a r t a r   o m   � v e r f � r i n g . o M � l k a t a l o g e n   i n n e h � l l e r   d e n   d e l v i s   � v e r f � r d a   f i l e n   ' % s ' ,   s o m   � r   s t � r r e   � n   k � l l f i l e n .   F i l e n   k o m m e r   a t t   t a s   b o r t . u * * V i l l   d u   l � g g a   t i l l   f i l e n   ' % s '   i   s l u t e t   a v   b e f i n t l i g   f i l ? * * 
 
 T r y c k   ' N e j '   f � r   a t t   � t e r u p p t a   f i l � v e r f � r i n g e n   i s t � l l e t . 4 % s 
   
 N y :             	 % s   b y t e s ,   % s 
 B e f i n t l i g :   	 % s   b y t e s ,   % s ' F i l e n   ' % s '   � r   s k r i v s k y d d a d .   S k r i v   � v e r ? � * * S k r i v   � v e r   l o k a l   f i l   ' % s ' ? * * M � l k a t a l o g e n   i n n e h � l l e r   r e d a n   f i l e n   ' % s ' . 
 V � l j   o m   d u   v i l l   s k r i v a   � v e r   f i l e n   e l l e r   h o p p a   � v e r   d e n n a   � v e r f � r i n g   o c h   b e h � l l a   b e f i n t l i g   f i l . � * * S k r i v   � v e r   f j � r r f i l   ' % s ' ? * * M � l k a t a l o g e n   i n n e h � l l e r   r e d a n   f i l e n   ' % s ' . 
 V � l j   o m   d u   v i l l   s k r i v a   � v e r   f i l e n   e l l e r   h o p p a   � v e r   d e n n a   � v e r f � r i n g   o c h   b e h � l l a   b e f i n t l i g   f i l .           � V � r d   k o m m u n i c e r a r   i n t e   m e r   � n   n � g r a   ' % d '   s e k u n d e r .   V � n t a r   f o r t f a r a n d e . . . 
 
 O B S :   O m   p r o b l e m e t   u p p r e p a s ,   p r o v a   a t t   s t � n g a   a v   ' O p t i m e r a   s t o r l e k e n   p �   a n s l u t n i n g s b u f f e r t ' .    & � t e r a n s l u t 
 N y t t   n a & m n      T u n n e l   f � r   % s  L � s e n o r d  L � s e n o r d   f � r   n y c k e l  S e r v e r p r o m p t  A n v � n d a r n a m n  A & n v � n d a r n a m n :  S e r v e r p r o m p t :   % s  N y t t   l � s e n o r d  S & v a r :    A n v � n d e r   T I S   a u t e n t i s e r i n g . % s $ A n v � n d e r   K r y p t o k o r t   a u t e n t i s e r i n g . % s 
 & L � s e n o r d : 0 A n v � n d e r   t a n g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % s  N & u v a r a n d e   l � s e n o r d :  & N y t t   l � s e n o r d  & B e k r � f t a   n y t t   l � s e n o r d :  A u t e n t i s e r a r   t u n n e l   g e n o m   % s  � v e r f � r   m e d   e t t   a n n a t   n a m n  & N y t t   n a m n : g* * S e r v e r n s   c e r t i f i k a t   � r   i n t e   k � n t .   D u   h a r   i n g e n   g a r a n t i   f � r   a t t   s e r v e r n   � r   d e n   d a t o r   s o m   d u   t r o r   a t t   d e   � r . * * 
 
 S e r v e r c e r t i f i k a t e t s   d e t a l j e r   f � l j e r : 
 
 % s 
 
 O m   d u   l i t a r   p �   c e r t i f i k a t e t ,   t r y c k   p �   ' J a ' .   F � r   a t t   a n s l u t a   u t a n   a t t   l a g r a   c e r t i f i k a t   t r y c k e r   d u   p �   ' N e j ' .   F � r   a t t   a v b r y t a   a n s l u t n i n g e n   t r y c k e r   p �   A v b r y t . 
 
 V i l l   d u   f o r t s � t t a   a n s l u t a   o c h   l a g r a   c e r t i f i k a t e t ? - -   O r g a n i s a t i o n :   % s 
 | -   P l a t s :   % s 
 | -   A n n a t :   % s 
  % s ,   % s c U t g i v a r e : 
 % s 
 � m n e : 
 % s 
 G i l t i g :   % s   -   % s 
 
 F i n g e r a v t r y c k : 
 -   S H A - 2 5 6 :   % s 
 -   S H A - 1 :   % s 
 
 S a m m a n f a t t n i n g :   % s $ & L � s e n o r d s f r a s   f � r   k l i e n t c e r t i f i k a t : " L � s e n o r d s f r a s   f � r   k l i e n t c e r t i f i k a t   H * * V i l l   d u   k o n v e r t e r a   d e n   p r i v a t a   n y c k e l f i l e n   % s   t i l l   P u T T Y - f o r m a t ? * * 
 
 % s * * � r   d u   s � k e r   p �   a t t   d u   v i l l   � v e r f � r a   f l e r a   f i l e r   t i l l   e n   e n d a   f i l   ' % s '   i   e n   k a t a l o g   ' % s ' ? * * 
 
 F i l e r   k o m m e r   a t t   s k r i v a s   � v e r . 
 
 O m   d u   v e r k l i g e n   v i l l   � v e r f � r a   a l l a   f i l e r   t i l l   e n   k a t a l o g   ' % s ' ,   b e h � l l a   d e r a s   n a m n ,   s e   t i l l   a t t   d u   a v s l u t a r   s � k v � g e n   m e d   e t t   s n e d s t r e c k .  n y c k e l b y t e s a l g o r i t m  v � r d n y c k e l t y p  � t k o m s t n y c k e l - I D  � & t k o m s t n y c k e l - I D :  H e m l i g   � t k o m s t n y c k e l  H e m l i g   � t k o m s t & n y c k e l : [ D i r e k t   d u b b l e r i n g   a v   m a p p a r   s t � d s   i n t e .   A n v � n d   e n   d u b b l e r i n g   v i a   e n   l o k a l   t i l l f � l l i g   k o p i a .  A n g e   m � l   f � r   t e m p o r � r   l a g r i n g . ) T i m e o u t ,   v � n t a r   p �   a t t   s e r v e r n   s k a   s v a r a .  P r o x y - a u t e n t i s e r i n g  P r o x y   & a n v � n d a r n a m n :  P r o x y   & l � s e n o r d : - A l l a   f i l e r   i   m � l k a t a l o g e n   k o m m e r   a t t   r a d e r a s ! P F o r t s � t t   a t t   a n s l u t a   t i l l   e n   o k � n d   s e r v e r   o c h   l � g g   t i l l   d e s s   v � r d n y c k e l   i   c a c h e ?    % s   ( p o r t   % d ) / V � r d n y c k e l n   � r   i n t e   c a c h a d   f � r   d e n   h � r   s e r v e r n : E D u   h a r   i n g e n   g a r a n t i   f � r   a t t   s e r v e r n   � r   d e n   d a t o r   d u   t r o r   a t t   d e n   � r . ' V a r n i n g      p o t e n t i e l l t   s � k e r h e t s i n t r � n g ! ' D e t t a   b e t y d e r   a t t   a n t i n g e n   % s   e l l e r   % s . , s e r v e r a d m i n i s t r a t � r e n   h a r   � n d r a t   v � r d n y c k e l n H a t t   d u   h a r   f a k t i s k t   a n s l u t i t   t i l l   e n   a n n a n   d a t o r   s o m   l � t s a s   v a r a   s e r v e r n   N y c k e l f i n g e r a v t r y c k e t   f � r   % s   � r : G V � r d n y c k e l n   m a t c h a r   i n t e   d e n   s o m   W i n S C P   h a r   c a c h a t   f � r   d e n   h � r   s e r v e r n : j O m   d u   l i t a r   p �   d e n   h � r   v � r d e n ,   v � l j   % s   f � r   a t t   l � g g a   t i l l   n y c k e l n   t i l l   W i n S C P s   c a c h e   o c h   f o r t s � t t   a n s l u t a .  & G o d k � n n X O m   d u   v i l l   f o r t s � t t a   a n s l u t a   b a r a   e n   g � n g   u t a n   a t t   l � g g a   t i l l   n y c k e l n   i   c a c h e n ,   v � l j   % s .  A n s l u t   & e n   g � n g I O m   d u   i n t e   l i t a r   p �   d e n   h � r   v � r d e n ,   v � l j   % s   f � r   a t t   a v b r y t a   a n s l u t n i n g e n . � O m   d u   f � r v � n t a d e   d i g   d e n   h � r   f � r � n d r i n g e n ,   l i t a r   p �   d e n   n y a   n y c k e l n   o c h   v i l l   f o r t s � t t a   a t t   a n s l u t a   t i l l   s e r v e r n ,   v � l j   a n t i n g e n   % s   f � r   a t t   u p p d a t e r a   c a c h e n   e l l e r   v � l j   % s   f � r   a t t   l � g g a   t i l l   d e n   n y a   n y c k e l n   t i l l   c a c h e n   s a m t i d i g t   s o m   d e n / d e   g a m l a   b e h � l l s . D O m   d u   v i l l   f o r t s � t t a   a n s l u t a   m e n   u t a n   a t t   u p p d a t e r a   c a c h e n ,   v � l j   % s . p O m   d u   v i l l   a v b r y t a   a n s l u t n i n g e n   h e l t ,   v � l j   % s   f � r   a t t   a v b r y t a .   A t t   v � l j a   % s   � r   d e t   E N D A   g a r a n t e r a d e   s � k r a   v a l e t . 7 D e n   h � r   s e r v e r n   p r e s e n t e r a d e   e n   c e r t i f i e r a d   v � r d n y c k e l : m s o m   s i g n e r a d e s   a v   e n   a n n a n   c e r t i f i k a t u t f � r d a r e   � n   d e n / d e   W i n S C P   � r   k o n f i g u r e r a d   a t t   l i t a   p �   f � r   d e n n a   s e r v e r . \ D e n   n y c k e l n   m a t c h a r   i n t e   h e l l e r   n y c k e l n   s o m   W i n S C P   t i d i g a r e   h a d e   c a c h a t   f � r   d e n   h � r   s e r v e r n . 6 e n   a n n a n   c e r t i f i k a t u t f � r d a r e   � r   v e r k s a m   i   d e t t a   o m r � d e b s o m   i n t e   m a t c h a r   d e n   c e r t i f i e r a d e   n y c k e l   s o m   W i n S C P   t i d i g a r e   h a d e   c a c h e l a g r a t   f � r   d e n   h � r   s e r v e r n . � ( A t t   l a g r a   d e n   h � r   c e r t i f i e r a d e   n y c k e l n   i   c a c h e n   k o m m e r   I N T E   a t t   g � r a   a t t   d e s s   c e r t i f i k a t u t f � r d a r e   k a n   l i t a s   p �   f � r   n � g o n   a n n a n   n y c k e l   e l l e r   v � r d . )  S � k e r h e t s v a r n i n g = V i l l   d u   a c c e p t e r a   r i s k e n   o c h   f o r t s � t t a   m e d   d e n   h � r   s e s s i o n e n ? \ D e   f � r s t a   % s   s o m   s t � d s   a v   s e r v e r n   � r   % s ,   v i l k e t   � r   u n d e r   d e n   k o n f i g u r e r a d e   v a r n i n g s t r � s k e l n . CD e n   % s   s o m   v a l t s   f � r   d e n   h � r   s e s s i o n e n   � r   % s ,   s o m   m e d   d e n   h � r   s e r v e r n   � r   s � r b a r   f � r   ' T e r r a p i n ' - a t t a c k e n   C V E - 2 0 2 3 - 4 8 7 9 5 ,   v i l k e t   p o t e n t i e l l t   t i l l � t e r   e n   a n g r i p a r e   a t t   � n d r a   d e n   k r y p t e r a d e   s e s s i o n e n . 
 
 U p p g r a d e r i n g ,   p a t c h n i n g   e l l e r   a t t   o m k o n f i g u r e r a   d e n n a   S S H - s e r v e r   � r   d e t   b � s t a   s � t t e t   a t t   u n d v i k a   d e n n a   s � r b a r h e t ,   o m   m � j l i g t . � D u   k a n   o c k s �   u n d v i k a   d e n n a   s � r b a r h e t   g e n o m   a t t   � v e r g e   d e n   h � r   s e s s i o n e n ,   f l y t t a   % s   t i l l   u n d e r   r a d e n   ' v a r n a   n e d a n '   i   W i n S C P : s   S S H - c h i f f e r k o n f i g u r a t i o n   ( s �   a t t   e n   a l g o r i t m   u t a n   s � r b a r h e t e n   k o m m e r   a t t   v � l j a s )   o c h   s t a r t a   e n   n y   s e s s i o n .          C O R E _ I N F O R M A T I O N  J a  N e j G V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 P r i v a t   n y c k e l f i l :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s  V e r s i o n   % s   ( % s ) > O p e r a t i o n e n   s l u t f � r d e s   f r a m g � n g s r i k t .   A n s l u t n i n g e n   a v s l u t a d e s .  S F T P - % d : S F T P   p r o t o k o l l e t s   v e r s i o n   t i l l � t e r   i n t e   n a m n b y t e   p �   f i l e r . ' S e r v e r n   s t � d e r   i n g a   u t � k n i n g a r   a v   S F T P . ( S e r v e r n   s t � d e r   f � l j a n d e   S F T P   u t � k n i n g a r :     
 L � & g g   t i l l  E n d a s t   n & y a r e  V i s a r   h j � l p . S t � n g e r   a l l a   s e s s i o n e r   o c h   a v s l u t a r   p r o g r a m m e t    A n s l u t e r   t i l l   s e r v e r  S t � n g e r   s e s s i o n e n 4 L i s t a r   a n s l u t n a   s e s s i o n e r   e l l e r   v � l j e r   a k t i v   s e s s i o n  V i s a r   a k t u e l l   f j � r r k a t a l o g  B y t e r   a k t u e l l   f j � r r k a t a l o g  V i s a r   i n n e h � l l e t   i   f j � r r k a t a l o g  V i s a r   a k t u e l l   l o k a l   k a t a l o g  B y t e r   a k t u e l l   l o k a l   k a t a l o g ! L i s t a r   i n n e h � l l e t   i   l o k a l   k a t a l o g  T a r   b o r t   f j � r r f i l  T a r   b o r t   f j � r r k a t a l o g $ F l y t t a r   e l l e r   b y t e r   n a m n   p �   f j � r r f i l   � n d r a r   r � t t i g h e t e r n a   p �   f j � r r f i l  S k a p a r   e n   s y m b o l i s k   f j � r r l � n k  S k a p a r   f j � r r k a t a l o g 3 L a d d a r   n e r   f i l   f r � n   f j � r r k a t a l o g   t i l l   l o k a l   k a t a l o g 3 L a d d a r   u p p   f i l   f r � n   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g - S � t t e r   e l l e r   v i s a r   v � r d e n   p �   s c r i p t a l t e r n a t i v , S y n k r o n i s e r a r   f j � r r k a t a l o g   m e d   l o k a l   k a t a l o g D K o n t i n u e r l i g t   � t e r s p e g l a   � n d r i n g a r   i   l o k a l   k a t a l o g   t i l l   f j � r r k a t a l o g  V � r d :      A k t i v   s e s s i o n :   [ % d ]   % s  S e s s i o n   ' % s '   a v s l u t a d .  L o k a l   ' % s '   % s   F j � r r   ' % s '  ' % s '   b o r t t a g e n 7 � v e r v a k a r   f � r � n d r i n g a r ,   t r y c k   C T R L - C   f � r   a t t   a v b r y t a . . .  & H o p p a   � v e r   a l l a  K � r   g o d t y c k l i g t   f j � r r k o m m a n d o  & T e x t  & B i n � r t   8 � v e r f � r i n g s t y p :   % s | B i n � r | T e x t | A u t o m a t i s k   ( % s ) | A u t o m a t i s k O F i l n a m n s f � r � n d r i n g :   % s | I n g e n   � n d r i n g | V e r s a l e r | G e m e n e r | F � r s t a   v e r s a l | G e m e n e r   8 . 3  S � t t   r � t t i g h e t e r :   % s  L � g g   t i l l   X   t i l l   k a t a l o g  B e v a r a   t i d s s t � m p e l    F i l m a s k :   % s  R e n s a   ' A r k i v '   a t t r i b u t  B y t   i n t e   u t   o g i l t i g a   t e c k e n    B e v a r a   i n t e   t i d s s t � m p e l  B e r � k n a   i n t e   � v e r f � r i n g s s t o r l e k   S t a n d a r d � v e r f � r i n g s i n s t � l l n i n g a r  V � r d n a m n :   % s  A n v � n d a r n a m n :   % s  F j � r r k a t a l o g :   % s    L o k a l   k a t a l o g :   % s $ S k a n n a r   ' % s '   e f t e r   u n d e r k a t a l o g e r . . . % � v e r v a k a r   � n d r i n g a r   i   % d   k a t a l o g e r . . .  � n d r i n g   i   ' % s '   u p p t � c k t .  F i l   ' % s '   � v e r f � r d .  F i l   ' % s '   b o r t t a g e n . U % s   k o n f i g u r e r a d   � v e r f � r i n g s i n s t � l l n i n g   k a n   i n t e   a n v � n d a s   i   a k t u e l l   k o n t e x t | N � g o n | A l l a    I g n o r e r a   r � t t i g h e t s f e l  A n v � n d e r   a n v � n d a r n a m n   " % s " . . A n v � n d e r   t a n g e n t b o r d s i n t e r a k t i v   a u t e n t i s e r i n g . % A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s " .  F e l a k t i g   l � s e n o r d .  � t k o m s t   n e k a d . 0 A u t e n t i s e r i n g   m e d   p u b l i k   n y c k e l   " % s "   f r � n   a g e n t . ( F � r s � k e r   m e d   p u b l i k   n y c k e l a u t e n t i s e r i n g . ' A u t e n t i s e r i n g   m e d   f � r i n s t � l l t   l � s e n o r d .  � p p n a r   t u n n e l . . .  A n s l u t n i n g   a v s l u t a d .    S � k e r   e f t e r   v � r d . . .  A n s l u t e r   t i l l   v � r d . . .  A u t e n t i s e r a r . . .  A u t e n t i s e r a d .  S t a r t a r   s e s s i o n e n . . .  L � s e r   f j � r r k a t a l o g . . .  S e s s i o n e n   s t a r t a d .  A n s l u t e r   g e n o m   t u n n e l . . .  S e r v e r   n e k a r   v � r   n y c k e l .  A d m i n i s t r a t i v t   f � r b j u d e n   ( % s ) .  A n s l u t n i n g   m i s s l y c k a d e s   ( % s ) . . N � t v e r k s f e l :   A n s l u t n i n g   t i l l   " % H O S T % "   n e k a d e s .   + N � t v e r k s f e l :   A n s l u t n i n g   � t e r s t � l l d   a v   p e e r . 5 N � t v e r k s f e l :   A n s l u t n i n g   t i l l   " % H O S T % "   g j o r d e   t i m e o u t . 2 V � r d :   % s 
 A n v � n d a r n a m n :   % s 
 � v e r f � r i n g s p r o t o k o l l :   % s 
 & � t e r u p p t a / S e r v e r n   s t � d e r   i n t e   n � g r a   e x t r a   F T P   e g e n s k a p e r . . S e r v e r n   s t � d e r   d e   h � r   e x t r a   F T P   e g e n s k a p e r n a :   # � v e r f � r i n g s h a s t i g h e t s g r � n s :   % u   k B / s  & K o p i e r a   n y c k e l 
 & U p p d a t e r a 
 & L � g g   t i l l  B e v a r a   e n d a s t   l � s n i n g 	 J � m f � r . . .  S y n k r o n i s e r a r . . .  I n g e t   a t t   s y n k r o n i s e r a . 
 O b e g r � n s a d  S S L / T L S   I m p l i c i t   k r y p t e r i n g      T L S / S S L   E x p l i c i t   k r y p t e r i n g  V i s a r   a r g u m e n t e n   s o m   m e d d e l a n d e  H � m t a r   a t t r i b u t   f � r   f j � r r f i l # V � r d e n s   f i n g e r a v t r y c k s n y c k e l   � r   % s . F V � x e l   - f i l e m a s k   � s i d o s � t t e r   f � r � l d r a d e   i n k l u d e r a / e x k l u d e r a   a l t e r n a t i v .  B a r a   & n y a   o c h   � n d r a d e   f i l e r � S e r v e r n   a v v i s a d e   S F T P - a n s l u t n i n g ,   m e n   d e n   l y s s n a r   p �   F T P - a n s l u t n i n g a r . 
 
 V i l l   d u   a n v � n d a   F T P - p r o t o k o l l e t   i s t � l l e t   f � r   S F T P ?   F � r e d r a r   a t t   a n v � n d a   k r y p t e r i n g . ` � p p n a   s e s s i o n   m e d   k o m m a n d o r a d s p a r a m e t e r   i   s k r i p t   � r   f � r � l d r a d .   A n v � n d   ' o p e n ' - k o m m a n d o t   i s t � l l e t . L V A R N I N G !   A t t   g e   u p p   s � k e r h e t e n   o c h   a c c e p t e r a   n � g o n   n y c k e l   s o m   k o n f i g u r e r a t s ! P V A R N I N G !   A t t   g e   u p p   s � k e r h e t e n   o c h   a c c e p t e r a   n � g o t   c e r t i f i k a t   s o m   k o n f i g u r e r a t s !  N y   l o k a l   f i l   % s  N y   f j � r r f i l   % s $ L o k a l   f i l   % s   � r   n y a r e   � r   f j � r r f i l   % s $ F j � r r f i l   % s   � r   n y a r e   � n   l o k a l   f i l   % s  � v e r g e   f j � r r f i l   % s  � v e r g e   l o k a l   f i l   % s  S k i l l n a d e r   h i t t a d e :  T a   b o r t   E O F - t e c k e n  T a   b o r t   B O M [ A n v � n d a   k o n f i g u r e r a d e   � v e r f � r i n g s i n s t � l l n i n g a r   s o m   s k i l j e r   s i g   f r � n   f a b r i k s i n s t � l l n i n g a r n a . \ A n v � n d a   k o n f i g u r e r a d e   s y n k r o n i s e r i n g s a l t e r n a t i v   s o m   s k i l j e r   s i g   f r � n   f a b r i k s i n s t � l l n i n g a r n a .    V e r s i o n  U t v e c k l i n g s v e r s i o n  F e l s � k n i n g s v e r s i o n  -   D i s t r i b u e r a   I N T E ' S e r v e r n   s t � d e r   d e s s a   W e b D A V   u t � k n i n g a r :  E x k l u d e r a   & k a t a l o g e r " B e r � k n a r   k o n t r o l l s u m m a   a v   f j � r r f i l    L a d d a r   k l i e n t c e r t i f i k a t . . . < S e r v e r n   f r � g a r   e f t e r   a u t e n t i s e r i n g   m e d   e t t   k l i e n t c e r t i f i k a t .  L � s t  K � r b a r � S k r i p t   a n v � n d e r   i n t e   f r i s t � e n d e   p a r a m e t r a r .   P a r a m e t r a r n a   d u   h a r   a n g e t t   p �   k o m m a n d o r a d e n   k o m m e r   i n t e   a t t   a n v � n d a s .   D i n   k o m m a n d o r a d s y n t a x   � r   f � r m o d l i g e n   f e l . Z I   s k r i p t ,   b � r   d u   a n v � n d a   e n   - h o s t k e y   v � x e l   f � r   a t t   k o n f i g u r e r a   d e n   f � r v � n t a d e   v � r d n y c k e l n . Y I   s k r i p t   s k a   d u   i n t e   f � r l i t a   d i g   p �   s p a r a d e   w e b b p l a t s e r ,   a n v � n d a   d e t t a   k o m m a n d o   i s t � l l e t :  K o n f i g u r e r a   s e s s i o n s a l t e r n a t i v  A n s l u t    L a d d a   W i n S C P   . N E T   a s s e m b l e r  % s   ( i n k l u s i v e   k a t a l o g e r ) , F i l e n   m � s t e   v a r a   k o d a d   i   U T F - 8   e l l e r   U T F - 1 6 . 	 % s   o c h   % s  � n d r a r   l � s e n o r d .  & K l i s t r a   i n   n y c k e l  D u p l i c e r a r   f j � r r f i l e n    O k � n d   ) & K o p i e r a   n y c k e l f i n g e r a v t r y c k   t i l l   u r k l i p p . & K o p i e r a   c e r t i f i k a t   f i n g e r a v t r y c k   t i l l   u r k l i p p  K r y p t e r a   i n t e   n y a   f i l e r  E x k l u d e r a   d o l d a   f i l e r  E x k l u d e r a   t o m m a   k a t a l o g e r U * * P u b l i k   n y c k e l   " % s "   i n s t a l l e r a d e s . * * 
 
 D u   k a n   n u   l o g g a   i n   p �   s e r v e r n   m e d   n y c k e l p a r e t . l E v e n t u e l l a   f e l   b e h � r i g h e t e r   f � r   f i l e n   " % s "   o c h / e l l e r   d e s s   f � r � l d r a m a p p   u p p t � c k t e s .   V � n l i g e n   k o n t r o l l e r a   d e m . � n y s s | i d a g | i g � r | i   m o r g o n | e n   s e k u n d   s e d a n | % d   s e k u n d e r   s e d a n | e n   m i n u t   s e d a n | % d   m i n u t e r   s e d a n | e n   t i m m e   s e d a n | % d   t i m m a r   s e d a n | e n   d a g   s e d a n | % d   d a g a r   s e d a n | e n   v e c k a   s e d a n |   % d   v e c k o r   s e d a n | e n   m � n a d   s e d a n | % d   m � n a d e r   s e d a n | e t t   � r   s e d a n | % d   � r   s e d a n  % d   d a g a r 5 B l � d d r a   e f t e r   I N I - f i l   a t t   i m p o r t e r a   w e b b p l a t s e r   f r � n . - L � g g e r   t i l l   p u b l i k   n y c k e l r a d   t i l l   f i l e n   " % s " :  H � m t a r   a k t u e l l   " % s " - f i l . . . 0 " % s " - f i l e n   i n n e h � l l e r   r e d a n   e n   p u b l i k   n y c k e l r a d : 8 " % s " - f i l e n   i n n e h � l l e r   i n t e   d e n   p u b l i k a   n y c k e l r a d e n   � n n u .    S k a p a r   n y   " % s " - f i l . . .   L a d a r   u p p   u p p d a t e r a d   " % s " - f i l . . .                                                C O R E _ V A R I A B L E ( S S H   o c h   S C P   k o d e n   � r   b a s e r a d   p �   P u T T Y   % s   " C o p y r i g h t   �   1 9 9 7  2 0 2 5   S i m o n   T a t h a m 3 h t t p s : / / w w w . c h i a r k . g r e e n e n d . o r g . u k / ~ s g t a t h a m / p u t t y /  F T P - k o d   b a s e r a d   p �   F i l e Z i l l a    C o p y r i g h t   �   T i m   K o s s e    h t t p s : / / f i l e z i l l a - p r o j e c t . o r g / m D e n n a   p r o d u k t   i n n e h � l l e r   p r o g r a m v a r a   s o m   u t v e c k l a t s   a v   O p e n S S L   P r o j e c t   f � r   a n v � n d n i n g   i   O p e n S S L : s   v e r k t y g   % s . ' C o p y r i g h t   �   1 9 9 8  % s   T h e   O p e n S S L   P r o j e c t    h t t p s : / / o p e n s s l - l i b r a r y . o r g / + W e b D A V / H T T P - k o d   b a s e r a d   p �   n e o n b i b l i o t e k   % s  C o p y r i g h t   �   1 9 9 9  2 0 2 5   J o e   O r t o n  h t t p s : / / n o t r o j . g i t h u b . i o / n e o n /  e X p a t   l i b r a r y   % s    h t t p s : / / l i b e x p a t . g i t h u b . i o /               ? h t t p s : / / w w w . c h i a r k . g r e e n e n d . o r g . u k / ~ s g t a t h a m / p u t t y / l i c e n c e . h t m l            * *  $ $ $ S 3 - k o d   b a s e r a d   p �   l i b s 3 - b i b l i o t e k   % s  C o p y r i g h t   �   B r y a n   I s c h o  h t t p s : / / g i t h u b . c o m / b j i / l i b s 3 0 h t t p s : / / g i t h u b . c o m / b j i / l i b s 3 / b l o b / m a s t e r / L I C E N S E                               & F e l   v i d   h � m t n i n g   a v   f i l l i s t a   f � r   " % s " . g C e r t i f i k a t   u t f � r d a d e s   i n t e   f � r   d e n   h � r   s e r v e r n .   D u   k a n s k e   a n s l u t e r   t i l l   e n   s e r v e r   s o m   l � t s a s   v a r a   " % s " . " I n g e n   f i l   m a t c h a n d e   ' % s '   h i t t a d e s . 0 V i s s a   c e r t i f i k a t   i   c e r t i f i k a t k e d j a n   � r   o g i l t i g a .    C e r t i f i k a t e t   � r   g i l t i g t . ! W e b D A V - r e s u r s   f l y t t a d e   t i l l   ' % s ' .  F � r   m � n g a   o m d i r i g e r i n g a r .  O m d i r i g e r i n g s l o o p   u p p t � c k t .  O g i l t i g   U R L   " % s " . ! P r o x y - a u t e n t i s e r i n g   m i s s l y c k a d e s . 1 V � r d n y c k e l   m a t c h a r   i n t e   k o n f i g u r e r a d   n y c k e l   " % s " ! < D e t   a n g i v n a   n a m n e t   k a n   i n t e   t i l l d e l a s   s o m   � g a r e   t i l l   e n   f i l . I D e t   a n g i v n a   n a m n e t   k a n   i n t e   t i l l d e l a s   s o m   d e n   p r i m � r a   g r u p p e n   f � r   e n   f i l . g D e n   b e g � r d a   � t g � r d e n   k u n d e   i n t e   s l u t f � r a s   e f t e r s o m   d e t   a n g i v n a   b y t e - i n t e r v a l l s l � s e t   i n t e   h a r   b e v i l j a t s . 7 P r i v a t   n y c k e l f i l   ' % s '   f i n n s   i n t e   e l l e r   k a n   i n t e   � p p n a s . & K o n t r o l l s u m m s a l g o r i t m   ' % s '   s t � d s   i n t e .  % s   % s   h a r   i n t e   v e r i f i e r a t s !   V a n l i g a   o r s a k e r   f � r   F e l k o d   4   � r : 
 -   B y t a   n a m n   p �   e n   f i l   t i l l   e t t   r e d a n   e x i s t e r a n d e   n a m n . 
 -   S k a p a   e n   k a t a l o g   s o m   r e d a n   f i n n s . 
 -   F l y t t a   e n   f j � r r f i l   t i l l   e t t   a n n a t   f i l s y s t e m   ( H D D ) . 
 -   � v e r f � r a   e n   f i l   t i l l   e t t   f u l l s t � n d i g t   f i l s y s t e m   ( H D D ) . 
 -   � v e r s k r i d a   e n   a n v � n d a r e s   d i s k k v o t .  K a n   i n t e   � p p n a   c e r t i f i k a t   " % s " .    K a n   i n t e   l � s a   c e r t i f i k a t   " % s " .   F e l   v i d   a v k o d n i n g   a v   c e r t i f i k a t . % F e l   v i d   a v k o d n i n g   a v   c e r t i f i k a t   " % s " . c C e r t i f i k a t f i l e n   " % s "   i n n e h � l l e r   i n t e   e n   p u b l i k   n y c k e l   o c h   i n g e n   m o t s v a r a n d e   . c r t / . c e r - f i l   h i t t a d e s .  F e l   v i d   l � s n i n g   a v   f i l e n   ' % s ' . ! F e l   v i d   u p p l � s n i n g   a v   f i l e n   ' % s ' .  F i l e n   ' % s '   � r   i n t e   l � s t . ) F e l   v i d   s p a r a n d e   a v   n y c k e l   t i l l   f i l   " % s " . K N e o n   H T T P - b i b l i o t e k e t s   i n i t i a l i s e r i n g   m i s s l y c k a d e s ,   k a n   i n t e   � p p n a   s e s s i o n . � V � l j a   f i l e r   m e d   h j � l p   a v   e t t   s � k v � g s s l u t   m e d   s n e d s t r e c k   � r   t v e t y d i g .   T a   b o r t   s n e d s t r e c k e t   f � r   a t t   v � l j a   m a p p .   B i f o g a   *   m a s k   f � r   a t t   v � l j a   a l l a   f i l e r   i   m a p p e n . � N � r   d u   a n s l u t e r   m e d   h j � l p   a v   e n   I P - a d r e s s ,   � r   d e t   i n t e   m � j l i g t   a t t   k o n t r o l l e r a   o m   c e r t i f i k a t e t   u t f � r d a d e s   f � r   s e r v e r n .   A n v � n d   e t t   v � r d n a m n   i s t � l l e t   f � r   I P - a d r e s s e n . E F � r v � n t a d e   v � r d n y c k e l   h a r   i n t e   k o n f i g u r e r a t s ,   a n v � n d   - h o s t k e y   s w i t c h . * O m d i r i g e r a s   t i l l   e n   o k r y p t e r a d   w e b b a d r e s s .  M o t t o g   s v a r   % d   " % s "   f r � n   % s . 2 F i l e Z i l l a   w e b b p l a t s h a n t e r a r f i l   h i t t a d e s   i n t e   ( % s ) . @ I n g a   w e b b p l a t s e r   h i t t a d e s   i   F i l e Z i l l a   w e b b p l a t s h a n t e r a r f i l   ( % s ) . ' F i l e Z i l l a   w e b b p l a t s   " % s "   h i t t a d e s   i n t e . [ D u   k a n   i n t e   a n s l u t a   t i l l   e n   S F T P - s e r v e r   m e d   h j � l p   a v   e n   F T P - p r o t o k o l l .   V � l j   r � t t   p r o t o k o l l . - F e l   u p p s t o d   v i d   l o g g n i n g .   K a n   i n t e   f o r t s � t t a .  ' % s '   � r   i n t e   e n   g i l t i g   s t o r l e k . ( O p e n S S H   f i l e n   k n o w n _ h o s t s   h i t t a d e s   i n t e . % I n g a   v � r d n y c k l a r   f i n n s   i   k n o w n _ h o s t s . R U r k l i p p e t s   i n n e h � l l   s t � m m e r   i n t e   � v e r e n s   m e d   v � r d n y c k e l n   e l l e r   d e s s   f i n g e r a v t r y c k . 
 R e s u r s :   % s  Y t t e r l i g a r e   d e t a l j e r :   % s  E x t r a   d e t a l j e r :  � t k o m s t   n e k a d . / F i l e n   � r   i n t e   k r y p t e r a d   m e d   e n   k � n d   k r y p t e r i n g . � * * O g i l t i g   k r y p t e r i n g s n y c k e l . * * 
 
 K r y p t e r i n g s n y c k e l n   f � r   k r y p t e r i n g   % s   m � s t e   h a   % d   b y t e .   D e n   m � s t e   a n g e s   i   h e x a d e c i m a l   r e p r e s e n t a t i o n   ( d v s   % d   t e c k e n ) . ) S e r v e r   s k i c k a d e   e n   f i l   s o m   i n t e   b e g � r d e s . & D e t   g i c k   i n t e   a t t   l a g r a   n y   v � r d n y c k e l . [ N � r   d u   l a d d a r   u p p   s t r e a m a d   d a t a   k a n   e n d a s t   e n   k � l l a   a n g e s   o c h   m � l e t   m � s t e   a n g e   e t t   f i l n a m n .   # F e l   v i d   l � s n i n g   a v   i n m a t n i n g s s t r � m . 2 F e l   v i d   l � s n i n g   a v   A W S - k o n f i g u r a t i o n s p a r a m e t e r   % s . o K a n   i n t e   s k a p a   t e m p o r � r   k a t a l o g   ' % s ' .   D u   k a n   � n d r a   r o t k a t a l o g e n   f � r   l a g r i n g   a v   t e m p o r � r a   f i l e r   i   I n s t � l l n i n g a r . * O p e n S S H - k o n f i g u r a t i o n s f i l e n   h i t t a d e s   i n t e . N I n g a   v � r d d i r e k t i v   f � r   s p e c i f i k a   v � r d a r   h i t t a d e s   i   O p e n S S H - k o n f i g u r a t i o n s f i l e n . + F T P - s e r v e r n   r e t u r n e r a d e   o g i l t i g t   s v a r   ' % s ' . K S 3 - p r o f i l e n   " % s "   e x i s t e r a r   i n t e   e l l e r   i n n e h � l l e r   i n g a   r e l e v a n t a   a l t e r n a t i v . 6 C e r t i f i k a t f i l e n   " % s "   f i n n s   i n t e   e l l e r   k a n   i n t e   � p p n a s . - D e t   g i c k   i n t e   a t t   l a d d a   c e r t i f i k a t f i l e n   " % s " . " U n k n o w n   p u b l i c   k e y   a l g o r i t h m   " % s " . C C e r t i f i k a t e t   i   " % s "   m a t c h a r   i n t e   d e n   p u b l i k a   n y c k e l n   i   n y c k e l f i l e n . ? D e t   g � r   i n t e   a t t   k o m b i n e r a   c e r t i f i k a t   i   " % s "   m e d   p r i v a t   n y c k e l . 6 F i l e n   " % s "   � r   i n t e   e n   p u b l i k   n y c k e l   i   e t t   k � n t   f o r m a t . . F i l e n s   s t o r l e k   " % s "   � r   % s ,   m e n   % s   f � r v � n t a d e s . ) I n l o g g n i n g s u p p g i f t e r   s p e c i f i c e r a d e s   i n t e .  K a n   i n t e   a v k o d a   n y c k e l :   % s ! O g i l t i g   n y c k e l   ( i n g e n   n y c k e l t y p ) . 9 C A - n y c k e l n   k a n s k e   i n t e   � r   e t t   c e r t i f i k a t   ( t y p e n   � r   ' % s ' ) .  O g i l t i g   n y c k e l d a t a   f � r   ' % s ' .                   " F e l   v i d   a n t a g a n d e t   a v   r o l l e n   ' % s ' . ! O v � n t a t   s v a r   p �   A W S - b e g � r a n   ( % s ) . ! I n g a   w e b b p l a t s e r   h i t t a d e s   i   " % s " . � S e r v e r n   a n v � n d e r   e t t   p r o t o k o l l   s o m   i n t e   s t � d s .   D i n   W i n S C P - s e s s i o n   � r   k o n f i g u r e r a d   a t t   a n v � n d a   % s   v i a   % s .   D e n   k a n   k o n f i g u r e r a s   f � r   a t t   a n v � n d a   % s   v i a   % s .   U n d v i k   d o c k   a t t   a n v � n d a   g a m l a   o s � k r a   p r o t o k o l l   n � r   d e t   � r   m � j l i g t .    O p e n S S L - i n i t i e r i n g   m i s s l y c k a d e s ( I n g e n   p r i v a t   n y c k e l   h i t t a d e s   i   f i l e n   % s .                                                       	 W I N _ E R R O R   Q % s 
   
 V a r n i n g :   A t t   a v b r y t a   d e n   h � r   o p e r a t i o n e n   k o m m e r   a t t   s t � n g a   n e r   a n s l u t n i n g e n !          K a n   i n t e   s k a p a   g e n v � g . ) K a n   i n t e   s k r i v a   � v e r   s p e c i a l s e s s i o n   ' % s ' .  K a n   i n t e   u t f o r s k a   k a t a l o g   ' % s ' . + I n g e n   f i l l i s t a   f � r   � v e r f � r i n g   h a r   a n g i v i t s .  K a n   i n t e   s k a p a   k a t a l o g e n   ' % s ' .   ' K a n   i n t e   t a   b o r t   t e m p o r � r   k a t a l o g   ' % s ' . % K a n   i n t e   � p p n a   e l l e r   k � r a   f i l e n   ' % s ' .  K a n   i n t e   s t a r t a   e d i t o r   ' % s ' .   w K a n   i n t e   � p p n a   m o t s v a r a d e   k a t a l o g   i   m o t s a t t   p a n e l .   S y n k r o n i s e r i n g   a v   k a t a l o g b l � d d r i n g   m i s s l y c k a d e s .   D e n   h a r   s t � n g t s   a v .  K a n   i n t e   a v g � r a   g e n v � g   ' % s ' .   % ' % s '   � r   i n t e   g i l t i g t   p r o f i l p l a t s n a m n . 4 ' % s '   � r   i n t e   g i l t i g t   n a m n   f � r   e n   p r o f i l p l a t s k a t a l o g . 1 P r o f i l p l a t s k a t a l o g e n   m e d   n a m n e t   ' % s '   f i n n s   r e d a n . 5 B e s k r i v n i n g   p �   e g e t   k o m m a n d o   k a n   i n t e   i n n e h � l l a   ' % s ' . 1 E g e t   k o m m a n d o   m e d   b e s k r i v n i n g e n   ' % s '   f i n n s   r e d a n . D K a n   i n t e   f r � g a   a p p l i k a t i o n e n s   h e m s i d a   e f t e r   u p p d a t e r i n g s i n f o r m a t i o n . , F e l   u p p s t o d   v i d   s � k n i n g   e f t e r   u p p d a t e r i n g a r .         < K a n   i n t e   r e g i s t r e r a   p r o g r a m m e t   f � r   a t t   h a n t e r a   U R L - a d r e s s e r . 2 M u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . E S k a l   d r a - t i l l � g g e t   m u t e x   s l � p p t e s   i n t e   e n l i g t   d e t   k r � v d a   i n t e r v a l l e t . �* * W i n S C P   k u n d e   i n t e   i d e n t i f i e r a   k a t a l o g e n ,   s o m   f i l e n   s l � p p t e s   i . * *   A n t i n g e n   h a r   d u   i n t e   s l � p p t   f i l e n   i   e n   v a n l i g   k a t a l o g   ( t . e x .   U t f o r s k a r e n )   e l l e r   o m   d u   i n t e   h a r   s t a r t a t   o m   d a t o r n   � n n u   e f t e r   i n s t a l l a t i o n e n   a v   s k a l t i l l � g g e t   d r a   &   s l � p p .   
 
 A l t e r n a t i v t   k a n   d u   v � x l a   t i l l   k o m p a t i b e l   d r a   &   s l � p p l � g e   ( f r � n   i n s t � l l n i n g s f � n s t r e t ) ,   s o m   a n v � n d e r   t e m p o r � r a   k a t a l o g e r   f � r   n e d l a d d n i n g a r .   D e t   g � r   a t t   d u   s l � p p a   f i l e r   t i l l   a l l a   d e s t i n a t i o n e r . K F i l e n   ' % s '   i n n e h � l l e r   i n t e   n � g o n   � v e r s � t t n i n g   f � r   d e n   h � r   p r o d u k t v e r s i o n e n . 5 F i l e n   ' % s '   i n n e h � l l e r   � v e r s � t t n i n g   f � r   % s   v e r s i o n   % s .   8 G S S A P I / S S P I   m e d   K e r b e r o s   s t � d s   i n t e   p �   d e t   h � r   s y s t e m e t . ' F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r . 8 F e l   u p p s t o d   v i d   b e v a k n i n g   a v   � n d r i n g a r   i   k a t a l o g e n   ' % s ' .   6 F e l   u p p s t o d   v i d   b e v a k n i n g e n   a v   � n d r i n g a r   i   f i l e n   ' % s ' . � * * K a n   i n t e   � v e r f � r a   d e n   r e d i g e r a d e   f i l e n   ' % s ' * * 
 
 S e s s i o n e n   ' % s '   h a r   r e d a n   s t � n g t s . 
 
 � p p n a   e n   n y   s e s s i o n   p �   s a m m a   w e b b p l a t s   o c h   f � r s � k   s p a r a   f i l e n   i g e n . I D e t   f i n n s   r e d a n   f � r   m � n g a   f i l e r   � p p n a d e .   V a r   g o d   s t � n g   n � g r a   f i l e r   f � r s t .   R % s   V a r   v � n l i g   t a   b o r t   f i l e n .   A n n a r s   k o m m e r   i n t e   a p p l i k a t i o n e n   a t t   f u n g e r a   k o r r e k t .   �W i n S C P   k u n d e   i n t e   a v g � r a   v i l k e t   p r o g r a m   s o m   s k a   s t a r t a s   f � r   a t t   � p p n a   f i l e n .   W i n S C P   k a n   i n t e   b e v a k a   � n d r i n g a r   i   f i l e n ,   s �   d e n   v i l l   i n t e   l a d d a s   u p p . 
   
 E n   m � j l i g   o r s a k   t i l l   p r o b l e m e t   � r   a t t   f i l e n   r e d a n   h a r   � p p n a t s   a v   e t t   a n n a t   p r o g r a m   s o m   k � r s . 
   
 O m   d u   v i l l   a n v � n d a   p r o g r a m m e t   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r . 
   
 N o t e r a   a t t   f i l e n   l i g g e r   k v a r   i   d e n   t e m p o r � r a   k a t a l o g e n . � N � g r a   a v   d e   t e m p o r � r a   k a t a l o g e r n a   k u n d e   i n t e   t a s   b o r t .   O m   f i l e r   f i n n s   l a g r a d e   d � r   s o m   f o r t f a r a n d e   � r   � p p n a ,   s t � n g   d e s s a   o c h   p r o v a   i g e n . � F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o ,   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   e n a   p a n e l e n ,   f � r   a t t   k � r a   k o m m a n d o t   p �   d e   v a l d a   f i l e r n a   i   m o t s a t t   p a n e l .   A l t e r n a t i v t   k a n   s a m m a   a n t a l   f i l e r   m a r k e r a s   i   b � d a   p a n e l e r n a   f � r   a t t   k � r a   k o m m a n d o t   p �   m a t c h a n d e   p a r   a v   f i l e r . W F � r   a t t   a n v � n d a   v a l t   e g e t   k o m m a n d o t   f � r   b a r a   e n   f i l   v a r a   m a r k e r a d   i   d e n   l o k a l a   p a n e l e n .   � N � g r a   a v   d e   v a l d a   f j � r r f i l e r n a   l a d d a d e s   i n t e   n e r .   D e t   v a l d a   e g n a   k o m m a n d o t   m � s t e   k � r a s   p �   m a t c h a n d e   p a r   a v   f i l e r ,   v i l k e t   d � r f � r   i n t e   � r   m � j l i g t . $ K a n   i n t e   i n i t i a l i s e r a   e x t e r n   k o n s o l .   N K a n   i n t e   � p p n a   m a p p n i n g s o b j e k t   f � r   a t t   s t a r t a   k o m m u n i k a t i o n   m e d   e x t e r n   k o n s o l . ; T i m e o u t   v � n t a r   p �   e x t e r n   k o n s o l   f � r   a t t   s l u t f � r a   k o m m a n d o t . 4 I n k o m p a t i b e l t   p r o t o k o l l v e r s i o n   f � r   e x t e r n   k o n s o l   % d . D F e l   u p p s t o d   n � r   s � k v � g   ' % s '   l a d e s   t i l l   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) . H F e l   u p p s t o d   n � r   s � k v � g   ' % s '   t o g s   b o r t   f r � n   m i l j � v a r i a b e l   p a t h ( % % P A T H % % ) .   [ F i l e n   ' % s '   � r   r e d a n   � p p n a d   i   e n   e x t e r n   e d i t o r   ( a p p l i k a t i o n )   e l l e r   h � l l e r   p �   a t t   l a d d a s   u p p . 8 D u   h a r   i n t e   a n g i v i t   n � g o n   a u t o m a t i s k t   v a l   a v   m a s k r e g l e r . D F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   m e d   b e s k r i v n i n g   ' % s '   f i n n s   r e d a n . x * * A n p a s s a t   k o m m a n d o   ' % s '   k a n   i n t e   k � r a s   j u s t   n u . * *   D u   k a n   b e h � v a   v � l j a   f i l e r   f � r   k o m m a n d o t   e l l e r   � p p n a   e n   s e s s i o n   f � r s t . A K a n   i n t e   l a d d a   o m   f i l e n   ' % s ' ,   s e s s i o n e n   ' % s '   h a r   r e d a n   a v s l u t a t s .         L � s e n o r d e t   k a n   i n t e   d e k r y p t e r a s . 3 D u   h a r   i n t e   a n g e t t   k o r r e k t   n u v a r a n d e   h u v u d l � s e n o r d . 0 N y a   o c h   u p p r e p a d e   h u v u d l � s e n o r d e t   � r   i n t e   s a m m a .   F E x t e r n   k o n s o l u t d a t a   d i r i g e r a s   t i l l   p i p e .   S e   t i l l   a t t   p i p e n   l � s e s   f r � n . ) ' % s '   � r   a r b e t s y t a ,   i n t e   w e b b p l a t s k a t a l o g . ) ' % s '   � r   w e b b p l a t s k a t a l o g ,   i n t e   a r b e t s y t a .   A K a n   i n t e   l � g g a   t i l l   s � k v � g   t i l l   % P A T H % ,   % P A T H %   � r   r e d a n   f � r   l � n g . 
 S t a c k s p � r :     A I n g a   w e b b p l a t s e r   h i t t a d e s   i   % s   r e g i s t e r n y c k e l   f � r   w e b b p l a t s   ( % s ) .   I n g e n   w e b b p l a t s m a s k   s p e c i f i c e r a d * I n g a   w e b b p l a t s i n s t � l l n i n g a r   s p e c i f i c e r a d e .  I n t e   � n d r a d  � n d r a d . H i t t a d e   % d   w e b b p l a t s e r ,   � n d r a d e   % d   w e b b p l a t s e r ! D u   m � s t e   a n g e   i n g � e n d e   n y c k e l f i l .  I n g e n   � t g � r d   a n g i v e n . " R e d i g e r a   S S H - 1   n y c k l a r   s t � d s   i n t e .  L � s e n f r a s e r n a   m a t c h a r   i n t e . ! D u   m � s t e   a n g e   u t g � e n d e   n y c k e l f i l . 4 F e l   v i d   h � m t n i n g   a v   u p p d a t e r i n g .   F � r s � k   i g e n   s e n a r e . E D e n   n e d l a d d a d e   u p p d a t e r i n g   k u n d e   i n t e   v e r i f i e r a s .   F � r s � k   i g e n   s e n a r e . C D i n   e - p o s t a d r e s s   h a r   i n t e   b e h � r i g h e t   f � r   a u t o m a t i s k a   u p p d a t e r i n g a r . F D i n   e - p o s t a d r e s s   b e h � r i g h e t   f � r   a u t o m a t i s k a   u p p d a t e r i n g a r   h a r   u p p h � r t . ^ D i n   e - p o s t a d r e s s   b l o c k e r a d e s   t i l l   a u t o m a t i s k a   u p p d a t e r i n g a r   p �   g r u n d   a v   � v e r d r i v e n   a n v � n d n i n g . � F � r   a t t   a k t i v e r a   a u t o m a t i s k a   u p p d a t e r i n g a r   f � r   d i n   e - p o s t a d r e s s ,   v � n l i g e n   f y l l   i   e t t   d o n a t i o n s f o r m u l � r   ( i n k l u s i v e   d i n   p o s t a d r e s s ) . 
 
 D u   h i t t a r   e n   l � n k   t i l l   f o r m u l � r e t   i   e t t   k v i t t o   s o m   d u   h a r   f � t t   e f t e r   d i n   d o n a t i o n . U D i n   d o n a t i o n   � r   u n d e r   d e n   g r � n s   s o m   k r � v s   f � r   a t t   a k t i v e r a   a u t o m a t i s k a   u p p d a t e r i n g a r . 
 I n g a   t i p s . & K o n v e r t e r a   p u b l i k a   n y c k l a r   s t � d s   i n t e .   / S � k e r   s e s s i o n   ( S S H   e l l e r   T L S / S S L )   i n t e   a n g i v e n .  U t � k n i n g e n   k r � v e r   % s . / O g i l t i g t   v � r d e   " % s "   f � r   u t � k n i n g s d i r e k t i v e t   % s . * S a k n a r   o b l i g a t o r i s k t   u t � k n i n g s d i r e k t i v   % s . " I n g e n   u t � k n i n g   f i n n s   i   d o k u m e n t e t . , D e t   f i n n s   r e d a n   e n   u t � k n i n g   m e d   n a m n e t   " % s " .   U t � k n i n g e n   � r   r e d a n   i n s t a l l e r a d . + F e l   v i d   i n l � s n i n g   a v   e n   u t � k n i n g   f r � n   " % s " . i * * I n g e n   s e s s i o n   � r   � p p e n * * 
 D e t   v a l d a   k o m m a n d o t   h a r   p l a t s s p e c i f i k a   a l t e r n a t i v ,   m e n   i n g e n   s e s s i o n   � r   � p p e n . (* * W i n S C P   k u n d e   i n t e   u p p t � c k a   e n   m a p p   d � r   d e   s l � p p t a   f i l e r n a   s l � p p t e s . * *   I   s t a n d a r d l � g e t   f � r   D r a   o c h   s l � p p   t i l l � t e r   W i n S C P   a t t   e n d a s t   f i l e r   s l � p p s   t i l l   l o k a l a   e n h e t e r   o c h   m a p p a d e   n � t v e r k s e n h e t e r . 
 
 D u   k a n   t i l l � t a   a t t   f i l e r   s l � p p s   t i l l   a n d r a   m � l   i   i n s t � l l n i n g a r .   T r y c k   p �   H j � l p - k n a p p e n   f � r   d e t a l j e r . " F e l   v i d   u p p d a t e r i n g   a v   s n a b b l i s t a .  F � r   m � n g a   p a r a m e t e r a r . ( S � k   i   i n k o r g e n   % s   e f t e r   " % s "   m e d d e l a n d e . ( I d e n t i t e t / n y c k e l f i l   s p e c i f i c e r a d e s   i n t e .  N y c k l a r   m � s t e   v a r a   u n i k a . ' T e c k n e t   " % s "   � r   i n t e   t i l l � t e t   i   t a g g a r .            W I N _ C O N F I R M A T I O N . S e s s i o n   m e d   n a m n   ' % s '   f i n n s   r e d a n .   S k r i v   � v e r ? ! K a t a l o g e n   ' % s '   f i n n s   i n t e .   S k a p a ?   � * * A v b r y t   f i l � v e r f � r i n g ? * * 
   
 O p e r a t i o n e n   k a n   i n t e   a v b r y t a s   i   m i t t e n   a v   f i l � v e r f � r i n g . 
 T r y c k   ' J a '   f � r   a t t   a v b r y t a   f i l � v e r f � r i n g   o c h   s t � n g a   a n s l u t n i n g e n . 
 T r y c k   ' N e j '   F � r   a t t   a v s l u t a   a k t u e l l   f i l � v e r f � r i n g . 
 T r y c k   ' A v b r y t '   f � r   a t t   f o r t s � t t a   o p e r a t i o n e n . . � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   f i l e n   ' % s ' ? 7 � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   d e   % d   v a l d a   f i l e r n a ? / A v s l u t a   s e s s i o n e n   ' % s '   o c h   s t � n g   a p p l i k a t i o n e n ?  F r � g a   m i & g   a l d r i g   i g e n 9F � r   l i t e   l e d i g t   u t r y m m e   p �   t e m p o r � r   e n h e t ! 
 
 N � r   f i l e r   d r a s   f r � n   e n   f j � r r k a t a l o g ,   l a d d a s   f i l e r n a   f � r s t   n e r   t i l l   e n   t e m p o r � r   k a t a l o g   ' % s ' .   D e t   � r   % s   l e d i g t   p �   e n h e t e n .   T o t a l   s t o r l e k   f � r   d e   v a l d a   f i l e r n a   � r   % s . 
 
 O B S :   T e m p o r � r   k a t a l o g e n   k a n   � n d r a s   i   I n s t � l l n i n g s f � n s t r e t . 
 
 V i l l   d u   f o r t s � t t a   m e d   a t t   l a d d a   n e r   f i l e r n a ?   ( L � g g   t i l l   k a t a l o g e n   ' % s '   t i l l   b o k m � r k e n ?     - S k a p a   g e n v � g   p �   s k r i v b o r d e t   f � r   s e s s i o n   ' % s ' ? 2 A n v � n d   a k t u e l l a   s e s s i o n s i n t � l l n i n g a r   s o m   s t a n d a r d ?  & H o p p a   � v e r # F i l e n   h a r   � n d r a t s .   S p a r a   � n d r i n g a r ? 9 S k a p a   u t f o r s k a r e n s   ' S k i c k a   t i l l ' - g e n v � g   f � r   s e s s i o n   ' % s ' ?  S k a p a   v a l d   i k o n / g e n v � g ? / A v s l u t a   a l l a   s e s s i o n e r   o c h   s t � n g   a p p l i k a t i o n e n ?   T a   b o r t   v a l d   p r o f i l p l a t s k a t a l o g ?  & F � r e g � e n d e  & N � s t a   3 V i l l   d u   r e g i s t r e r a   W i n S C P   a t t   h a n t e r a   U R L - a d r e s s e r ? L V i l l   d u   r e n s a   u p p   d a t a   f r � n   d e n   h � r   d a t o r n   s o m   h a r   s k a p a t s   a v   a p p l i k a t i o n e n ? ! % s 
 
 V i l l   d u   s t � n g a   a p p l i k a t i o n e n ? G % % s 
 
 V i l l   d u   a v s l u t a   % d   � t e r s t � e n d e   s e s s i o n e r   o c h   s t � n g a   a p p l i k a t i o n e n ? � * * D e t   f i n n s   f o r t f a r a n d e   n � g r a   � v e r f � r i n g a r   i   b a k g r u n d s k � n .   V i l l   d u   k o p p l a   n e r   i a l l a f a l l ? * * 
 
 V a r n i n g :   O m   d u   t r y c k e r   p �   ' O K '   k o m m e r   a l l a   � v e r f � r i n g a r   a t t   a v s l u t a s   o m e d e l b a r t . * * V i l l   d u   � p p n a   s e p a r a t   s k a l s e s s i o n ? * * 
 
 N u v a r a n d e   s e s s i o n   % s   s t � d e r   i n t e   k o m m a n d o t   d u   b e g � r .   S e p a r a t   s k a l s e s s i o n   k a n   � p p n a s   f � r   a t t   b e a r b e t a   k o m m a n d o t . 
 
 O B S :   S e r v e r n   m � s t e   e r b j u d a   U n i x - l i k n a n d e   s k a l   o c h   s k a l e t   m � s t e   a n v � n d a   s a m m a   s � k v � g s s y n t a x   s o m   n u v a r a n d e   s e s s i o n   % s . � D e t   f i n n s   n � g r a   � p p n a   f i l e r .   V a r   v � n l i g   s t � n g   d e m   i n n a n   a p p l i k a t i o n e n   a v s l u t a s . 
   
 O B S :   O m   d e t t a   i n t e   u t f � r s ,   k a n   r e d i g e r a d e   f i l e r   l i g g a   k v a r   i   d e n   t e m p o r � r a   k a t a l o g e n . '* * V i l l   d u   t a   b o r t   t i d i g a r e   t i l l f � l l i g a   k a t a l o g e r ? * * 
 
 W i n S C P   h a r   h i t t a t   % d   t e m p o r � r a   k a t a l o g e r ,   s o m   f � r m o d l i g e n   h a r   s k a p a t s   t i d i g a r e .   D e s s a   k a t a l o g e r   k a n   i n n e h � l l a   f i l e r   s o m   t i d i g a r e   h a r   r e d i g e r a t s   e l l e r   l a d d a t s   n e r . 
 
 D u   k a n   o c k s �   � p p n a   k a t a l o g e r   f � r   a t t   s e   � v e r   i n n e h � l l e t   o c h   t a   b o r t   d e m   s j � l v .  & � p p n a # V i s a   i n t e   d e t   h � r   m e d d e l a n d e t   i & g e n   f * * V i l l   d u   s k a p a   s k r i v b o r d s i k o n   f � r   a l l a   a n v � n d a r e ? * * 
 
 D u   m � s t e   h a   a d m i n i s t r a t � r s r � t t i g h e t e r   f � r   d e t t a . U V i l l   d u   l � g g a   t i l l   a p p l i k a t i o n e n s   s � k v � g   ' % s '   t i l l   m i l j � v a r i a b e l n s   s � k v � g   ( % % P A T H % % ) ? �E d i t o r n   ( a p p l i k a t i o n )   s o m   s t a r t a d e s   f � r   a t t   � p p n a   f i l   ' % s '   a v s l u t a d e s   f � r   t i d i g t .   O m   d e n   i n t e   a v s l u t a d e s   a v   e r ,   k a n   d e t   b e r o   p �   a t t   d e n   e x t e r n a   e d i t o r   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g a r e   s t a r t a d e   i n s t a n s e r   a v   e d i t o r n   s k i c k a r   s e d a n   d e n   n y a   f i l e n   t i l l   b e f i n t l i g a   i n s t a n s e r   a v   e d i t o r n   o c h   a v s l u t a r   s i g   o m e d e l b a r t .   F � r   a t t   s t � d j a   d e n n a   t y p   a v   e d i t o r s ,   m � s t e   W i n S C P   a n p a s s a   s i t t   b e t e e n d e ,   i n t e   t a   b o r t   t e m p o r � r   f i l   n � r   p r o c e s s e n   a v s l u t a r ,   u t a n   a t t   b e h � l l a   d e n   s �   l � n g e   W i n S C P   � r   i g � n g .   B e t e e n d e t   k a n   s t � n g a s   a v   g e n o m   a t t   � n d r a   i n s t � l l n i n g a r   f � r   e d i t o r n   ' E x t e r n   e d i t o r   � p p n a r   v a r j e   f i l   i   e t t   s e p a r a t   f � n s t e r   ( p r o c e s s ) ' .   O m   d i n   e d i t o r   i n t e   � r   a v   d e t   h � r   s l a g e t ,   b o r t s e   f r � n   d e t t a   m e d d e l a n d e   o c h   l � t   f i l e n   t a s   b o r t   f r � n   d e n   t e m p o r � r a   k a t a l o g e n   n u . 
   
 V i l l   n i   t a   b o r t   d e n   � p p n a d e   f i l e n   n u ?   ( G e n o m   a t t   t r y c k a   p �   ' N e j '   k o m m e r   d u   a t t   m � j l i g g � r a   d e t   s � r s k i l d a   b e t e e n d e t   o c h   b e h � l l a   f i l e n   i   t e m p o r � r a   k a t a l o g e n . )   � * * V i l l   d u   g � r a   r i k t n i n g e n   d u   v a l t   t i l l   s t a n d a r d ? * * 
 
 D u   h a r   � s i d o s a t t   f � r v a l d   s y n k r o n i s e r i n g s r i k t n i n g .   S o m   s t a n d a r d   b e s t � m s   r i k t n i n g e n   a v   f i l p a n e l e n   s o m   v a r   a k t i v   i n n a n   i n n a n   d u   k � r d e   s y n k r o n i s e r i n g s f u n k t i o n e n . � * * V i l l   d u   f � r s t   u t f � r a   e n   f u l l s t � n d i g   s y n k r o n i s e r i n g   a v   f j � r r k a t a l o g e n ? * * 
 
 F u n k t i o n e n   ' H � l l   f j � r r k a t a l o g   u p p d a t e r a d '   f u n g e r a r   k o r r e k t   e n d a s t   o m   f j � r r k a t a l o g e n   � r   s y n k r o n i s e r a d   m e d   d e n   l o k a l a   i n n a n   d e n   s t a r t a r . 1 S � k e r   p �   a t t   d u   v i l l   t a   b o r t   s p a r a d   s e s s i o n   ' % s ' ? � F l e r   � n   % d   k a t a l o g e r   o c h   u n d e r k a t a l o g e r   h i t t a d e s .   B e v a k n i n g   a v   � n d r i n g a r   i   m � n g a   k a t a l o g e r   k a n   s i g n i f i k a n t   m i n s k a   p r e s t a n d a n   p �   d a t o r n . 
   
 V i l l   d u   s k a n n a   f l e r   k a t a l o g e r ,   u p p   t i l l   % d   k a t a l o g e r ? 	 % s   ( % d   s )   8 S � k e r   p �   a t t   d u   v i l l   f l y t t a   f i l   ' % s '   t i l l   p a p p e r s k o r g e n ? > S � k e r   p �   a t t   d u   v i l l   f l y t t a   % d   v a l d a   f i l e r   t i l l   p a p p e r s k o r g e n ? I F i l e n   h a r   � n d r a t s .   � n d r i n g a r   v i l l   f � r l o r a s ,   o m   f i l e n   l a d d a s   o m .   F o r t s � t t ?  K & o n f i g u r e r a . . . ^ * * V i l l   d u   f � r s � k a   s k a p a   k a t a l o g e n   ' % s ' ? * * 
 
 K a n   i n t e   � p p n a   m o t s v a r a n d e   k a t a l o g   i   m o t s a t t   p a n e l .  L � g g   t i l l   & d e l a d e   b o k m � r k e n s* * V i l l   d u   s k i c k a   m e d d e l a n d e t   t i l l   W i n S C P : s   w e b b p l a t s ? * * 
 
 D e t   f i n n s   i n g e n   h j � l p s i d a   a s s o c i e r a d   m e d   m e d d e l a n d e t .   W i n S C P   k a n   s � k a   p �   s i n   d o k u m e n t a t i o n s p l a t s   e f t e r   m e d d e l a n d e t e x t e n . 
 
 O B S :   W i n S C P   k o m m e r   a t t   s k i c k a   m e d d e l a n d e t   � v e r   e n   o s � k e r   a n s l u t n i n g .   K o n t r o l l e r a   a t t   m e d d e l a n d e t   i n t e   i n n e h � l l e r   n � g o n   d a t a   s o m   d u   v i l l   s k y d d a ,   t i l l   e x e m p e l   n a m n   p �   f i l e r ,   k o n t o n   e l l e r   v � r d a r . 9* * D i t t   l � s e n o r d   � r   f � r   e n k e l t   o c h   k a n   i n t e   g e   t i l l r � c k l i g t   s k y d d   m o t   a t t a c k e r   m e d   o r d l i s t a   e l l e r   b r u t e   f o r c e . 
 � r   d u   s � k e r   a t t   d u   v i l l   a n v � n d a   d e t ? * * 
 
 O B S :   b r a   l � s e n o r d   h a r   m i n s t   s e x   t e c k e n   o c h   i n n e h � l l e r   b � d e   g e m e n e r   o c h   v e r s a l e r ,   s i f f r o r   o c h   s p e c i a l t e c k e n ,   s �   s o m   a v g r � n s a r e ,   s y m b o l e r ,   b o k s t � v e r   m e d   a c c e n t ,   e t c . 9 S k a p a   g e n v � g   p �   s k r i v b o r d e t   t i l l   w e b b p l a t s k a t a l o g e n   ' % s ' ? 0 S k a p a   g e n v � g   p �   s k r i v b o r d e t   t i l l   a r b e t s y t a   ' % s ' ? E V i l l   d u   � t e r a n s l u t a   s e s s i o n   ' % s '   f � r   a t t   � v e r f � r a   r e d i g e r a d   f i l   ' % s ' ? K A v s l u t a   a l l a   s e s s i o n e r   o c h   s t � n g   a p p l i k a t i o n e n   u t a n   a t t   s p a r a   e n   a r b e t s y t a ? � * * V i l l   d u   a n v � n d a   % s   i s t � l l e t   f � r   i n t e r n a   s t a n d a r d e d i t o r ? * * 
 
 W i n S C P   h a r   u p p t � c k t   a t t   d u   h a r   d e n   a n p a s s a d e   t e x t e d i t o r n   ' % s '   a s s o c i e r a d   m e d   t e x t f i l e r . � * * D u   h a r   s p a r a t   s e s s i o n e r / w e b b p l a t s e r   i   % s . 
 
 V i l l   d u   i m p o r t e r a   d e m   t i l l   W i n S C P ? * * 
 
 ( D u   k a n   i m p o r t e r a   d e m   n � r   s o m   h e l s t   s e n a r e   i   d i a l o g r u t a n   L o g g a   i n ) | P u T T Y   S S h - k l i e n t | F i l e z i l l a   F T P - k l i e n t | % s   o c h   % s  * * � t e r s t � l l   k o n f i g u r a t i o n   f r � n   e n   s � k e r h e t s k o p i a ? * * 
 
 I m p o r t   a v   k o n f i g u r a t i o n   k o m m e r   a t t   s k r i v a   � v e r   a l l a   d i n a   i n s t � l l n i n g a r   o c h   w e b b p l a t s e r .   W i n S C P   k o m m e r   a t t   s t a r t a s   o m   m e d   d e n   n y a   k o n f i g u r a t i o n e n .   � v e r v � g   a t t   s p a r a   d i t t   a r b e t e   o c h   s k a p a   e n   s � k e r h e t s k o p i a   a v   d i n   n u v a r a n d e   k o n f i g u r a t i o n .  & A l l a  J & a   t i l l   a l l a  R a & p p o r t e r a � D e t   f i n n s   a n d r a   i n s t a n s e r   a v   W i n S C P   i g � n g . 
 
 S t � l l a   i n   e l l e r   r e n s a   h u v u d l � s e n o r d e t ,   m e d a n   e n   a n n a n   i n s t a n s   a v   W i n S C P   � r   i g � n g ,   k a n   o r s a k a   f � r l u s t   a v   d i n a   l a g r a d e   l � s e n o r d . 
 
 V � n l i g e n   a v s l u t a   a n d r a   i n s t a n s e r   a v   W i n S C P   i n n a n   d u   f o r t s � t t e r . � V i l l   d u   b i f o g a   r e d i g e r a d   f i l   ' % s '   t i l l   s e s s i o n   ' % s ' ? * * 
 
 O r i g i n a l   s e s s i o n e n   s o m   a n v � n d e s   f � r   a t t   l a d d a   n e r   f i l e n   ' % s '   t i l l   e d i t o r n   h a r   r e d a n   s t � n g t s . @ V i l l   d u   a v r e g i s t r e r a   W i n S C P   f r � n   h a n t e r i n g   a v   a l l a   U R L - a d r e s s e r ? * * F � r s � k   a t t   � p p n a   s t o r   f i l ? * * 
 
 F i l e n   d u   f � r s � k e r   � p p n a   i   e n   i n t e r n   e d i t o r   � r   f � r   s t o r   ( % s ) .   W i n S C P   i n t e r n   e d i t o r   � r   i n t e   a v s e d d   f � r   r e d i g e r i n g   a v   s t o r a   f i l e r .   � v e r v � g   a t t   a n v � n d a   e n   e x t e r n   e d i t o r   s o m   k a n   r e d i g e r a   s t o r a   f i l e r . 
 
 D u   k a n   f � r s � k a   � p p n a   f i l e n   � n d � ,   m e n   W i n S C P   k a n   m i s s l y c k a s .  S t � n g X U t � k n i n g e n   k o m m e r   i n t e   f r � n   e n   b e t r o d d   k � l l a .   � r   d u   s � k e r   p �   a t t   d u   v i l l   i n s t a l l e r a   d e n ? � * * A n v � n d e r   d e n   s e n a s t e   k o m p a t i b l a   o c h   b e t r o d d a   v e r s i o n   a v   u t � k n i n g e n . * * 
 
 D e n   s e n a s t e   v e r s i o n e n   a v   u t � k n i n g e n   h a r   a n t i n g e n   i n t e   g r a n s k a t s   e l l e r   � r   i n t e   k o m p a t i b e l   m e d   d e n   h � r   v e r s i o n e n   a v   W i n S C P . [* * V i l l   d u   s k r i v a   � v e r   e n   b e f i n t l i g   I N I - f i l   ' % s ' ? * * 
 
 V � l j   ' S k r i v   � v e r '   f � r   a t t   s k r i v a   � v e r   d e n   v a l d a   I N I - f i l e n   m e d   d e n   a k t u e l l a   k o n f i g u r a t i o n e n . 
 
 V � l j   ' A n v � n d '   f � r   a t t   s t a r t a   o m   W i n S C P   m e d   e n   k o n f i g u r a t i o n   l a d d a d   f r � n   d e n   v a l d a   I N I - f i l e n .   D i n   n u v a r a n d e   k o n f i g u r a t i o n   k o m m e r   a t t   b e v a r a s   o c h   d u   k a n   � t e r g �   t i l l   d e n ,   o m   d e t   b e h � v s . | & S k r i v   � v e r | & A n v � n d =* * V i l l   d u   s k r i v a   � v e r   e n   s k r i v s k y d d a d   I N I - f i l   ' % s '   f � r   a t t   s p a r a   d i n   n u v a r a n d e   k o n f i g u r a t i o n ? * * D e n   h � r   f r � g a n   b l i r   i f r � g a s a t t   n � r   d u   h � l l e r   n e d   S h i f t - t a n g e n t e n   m e d a n   W i n S C P   s t � n g s   o c h   d i n   I N I - f i l   � r   s k r i v s k y d d a d .   N o r m a l t   s k r i v s   i n t e   I N I - f i l e r   � v e r   o c h   i n g a   � n d r i n g a r   i   k o n f i g u r a t i o n e n   g � r   f � r l o r a d e   n � r   W i n S C P   s t � n g s . K A v s l u t a   s e s s i o n e n   ' % s '   o c h   s t � n g   a p p l i k a t i o n e n   u t a n   a t t   s p a r a   e n   a r b e t s y t a ? - S t � n g   p r o g r a m m e t   u t a n   a t t   s p a r a   e n   a r b e t s y t a ? � * * V i l l   d u   v e r k l i g e n   � p p n a   e n   a n n a n   f l i k ? * * 
 D u   h a r   r e d a n   % d   f l i k a r   � p p n a .   � v e r v � g   a t t   s t � n g a   n � g r a   f l i k a r   f � r s t   f � r   a t t   f r i g � r a   r e s u r s e r   p �   d i n   d a t o r . M F j � r r f i l e n   h a r   � n d r a t s   m e d a n   d u   r e d i g e r a d e   d e n .   V i l l   d u   s k r i v a   � v e r   d e n   � n d � ?                      W I N _ I N F O R M A T I O N    I n g a   s k i l l n a d e r   h i t t a d e s .  � p p n a r   s e s s i o n   ' % s ' 
 % s ' V � n t a r   p �   a t t   d o k u m e n t e t   s k a   s t � n g a s . . .  % s   ( � v e r f � r   m e d   % s )  % s   ( f � r   � v e r f � r i n g )  L o k a l :   % s 
 F j � r r :   % s  & T o u c h  & K � r     1 % d   f e l   u p p s t o d   v i d   s e n a s t e   o p e r a t i o n e n .   V i s a   d e m ?  F e l   % d   a v   % d : 
 % s  D u   h a r   d e n   s e n a s t e   v e r s i o n e n .  N y   v e r s i o n   % s   h a r   s l � p p t s .  P a r a m e t e r v � r d e :  ' % s '   k o m m a n d o p a r a m e t r a r                      U R L :   P r o t o k o l l e t   % s  A n s l u t e r . . .  F r � g a  F e l  P r o m p t 	 V � n t a r . . .  T a & r / G Z i p . . .  & A r k i v n a m n :  & U n T a r / G Z i p . . .  P a c k a   & u p p   t i l l   k a t a l o g :    & G r e p . . .  & S � k   e f t e r   m � n s t e r :  % d   L � s e r   k a t a l o g  L i s t n i n g . . .    & U p p g r a d e r a   ; F � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s '   v a l d e s   a u t o m a t i s k t . 4 � t e r g �   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g   ' % s ' . + � t e r g �   t i l l   s t a n d a r d � v e r f � r i n g s i n s t � l l n i n g .  R e g e l   f � r   a u t o m a t i s k t   v a l : 
 % s    A d   H o c  P a u s a  & I n t e r n   e d i t o r �A p p l i k a t i o n   s t a r t a d   f � r   a t t   � p p n a   f i l   ' % s '   s t � n g d e s   f � r   t i d i g t .   O m   d e n   i n t e   s t � n g d e s   a v   d i g ,   d e   k a n   b e r o   p �   a t t   a p p l i k a t i o n e n   � p p n a r   f l e r a   f i l e r   i   e t t   f � n s t e r   ( p r o c e s s ) .   Y t t e r l i g a r e   s t a r t a d e   i n s t a n s e r   a v   a p p l i k a t i o n e n   s k i c k a r   d �   d e n   n y a   f i l e n   t i l l   b e f i n t l i g   a p p l i k a t i o n   o c h   s t � n g s   o m e d e l b a r t .   W i n S C P   k a n   s t � d j a   s � d a n a   a p p l i k a t i o n e r   e n d a s t   s o m   e x t e r n   e d i t o r . 
   
 O m   d u   v i l l   a n v � n d a   a p p l i k a t i o n e n   f � r   a t t   � p p n a   f i l e r   f r � n   W i n S C P ,   � v e r v � g a   a t t   k o n f i g u r e r a   d e n   s o m   e n   e x t e r n   e d i t o r .     = R e d i g e r a   ( e x t e r n ) | R e d i g e r a   v a l d a   f i l e r   m e d   e x t e r n   e d i t o r   ' % s ' � *   m a t c h a r   a l l a   a n t a l   t e c k e n . 
 ?   m a t c h a r   e x a k t   e t t   t e c k e n . 
 [ a b c ]   m a t c h a r   e t t   t e c k e n   f r � n   u p p s � t t n i n g e n . 
 [ a - z ]   m a t c h a r   e t t   t e c k e n   i   i n t e r v a l l e t . 
 E x e m p e l :   * . h t m l ;   p h o t o ? ? . p n g > M a s k   k a n   u t � k a s   m e d   s � k v � g s m a s k . 
 E x e m p e l :   * / p u b l i c _ h t m l / * . h t m l �M � n s t e r : 
 ! !   e x p a n d e r a r   t i l l   u t r o p s t e c k e n 
 !   e x p a n d e r a r   t i l l   f i l n a m n 
 ! &   e x p a n d e r a r   t i l l   l i s t a   m e d   v a l d a   f i l e r   ( c i t a t i o n s t e c k e n ,   m e l l a n s l a g s s e p a r e r a d ) 
 ! /   e x p a n d e r a r   t i l l   a k t u e l l   f j � r r s � k v � g 
 ! S   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s - U R L 
 ! @   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s v � r d n a m n 
 ! U   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s a n v � n d a r n a m n 
 ! P   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s l � s e n o r d 
 ! #   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   p o r t n u m m e r 
 ! N   e x p a n d e r a r   t i l l   a k t u e l l t   s e s s i o n s n a m n 
 ! ? p r o m p t [ \ ] ? d e f a u l t !   e x p a n d e r a r   t i l l   a n v � n d a r v a l t   v � r d e   m e d   g i v e n   p r o m p t   o c h   s t a n d a r d   ( a l t e r n a t i v t   \   u n d v i k e r   e s c a p e ) 
 ! ` c o m m a n d `   e x p a n d e r a r   t i l l   u t d a t a   a v   l o k a l t   k o m m a n d o 
   
 L o k a l t   k o m m a n d o m � n s t e r : 
 ! ^ !   e x p a n d e r a r   t i l l   f i l n a m n   f r � n   l o k a l   p a n e l 
   
 E x e m p e l : 
 g r e p   " ! ? M � n s t e r : ? ! "   ! & A A l l a   � v e r f � r i n g a r   i   b a k g r u n d e n   s l u t f � r d e s .   A n s l u t n i n g   a v s l u t a d e s .   L � s n i n g   a v   f j � r r k a t a l o g   a v b r � t s . ( S y n k r o n i s e r a d   b l � d d r i n g   s a t t e s   % s . | p � | a v ' V i s n i n g   a v   d o l d a   f i l e r   s a t t e s   % s . | p � | a v G A u t o m a t i s k   u p p d a t e r i n g   a v   f j � r r k a t a l o g   e f t e r   o p e r a t i o n   s a t t e s   % s . | p � | a v 1 � v e r f � r i n g   i   b a k g r u n d e n   k r � v e r   d i n   u p p m � r k s a m h e t .  � v e r f � r i n g s k � n   � r   t o m . Z ! Y   � r 
 ! M   m � n a d 
 ! D   d a g 
 ! T   t i d 
 ! P   p r o c e s s   i d 
 ! @   v � r d n a m n 
 ! S   s e s s i o n s n a m n 
 E x e m p e l : C : \ ! S ! T . l o g K P a s s i v t   l � g e   m � s t e   v a r a   a k t i v e r a d   n � r   F T P   a n s l u t n i n g   g e n o m   p r o x y   h a r   v a l t s . L U p p d a t e r i n g s k o n t r o l l   f � r   a p p l i k a t i o n e n   � r   t e m p o r � r t   a v s t � n g d .   F � r s � k   s e n a r e .  & G �   t i l l  V a d   � r   n y t t      O p e r a t i o n e n   s l u t f � r d e s  & P r i n t  & A s s o c i e r a d   a p p l i k a t i o n  P �  A v  A u t o S * * H u v u d l � s e n o r d e t   h a r   � n d r a t s . * * 
 
 D i n a   l a g r a d e   l � s e n o r d   � r   s � k r a d e   m e d   A E S - c h i f f e r .  H u v u d l � s e n o r d e t   h a r   � n d r a t s . S * * D u   h a r   t a g i t   b o r t   h u v u d l � s e n o r d e t . * * 
 
 D i n a   l a g r a d e   l � s e n o r d   � r   i n t e   s � k r a   l � n g r e .  H u v u d l � s e n o r d :      K o m m e r   a t t   k o n t r o l l e r a   i g e n :   % s  S e n a s t e   s e s s i o n e r Q M a s k e r   s k i l j s   � t   m e d   s e m i k o l o n   e l l e r   k o m m a .   
 P l a c e r a   u t e s l u t n a   m a s k e r   e f t e r   p i p e . , M a s k s l u t   m e d   s n e d s t r e c k   v � l j e r   u t   k a t a l o g e r .   � > s t o r l e k   m a t c h a r   f i l   s o m   � r   s t � r r e   � n   s t o r l e k 
 < s t o r l e k   m a t c h a r   f i l   m i n d r e   � n   s t o r l e k 
 > y y y y - m m - d d   m a t c h a r   f i l   s o m   � n d r a t s   e f t e r   d e t   d a t u m e t 
 < y y y y - m m - d d   m a t c h a r   f i l   s o m   � n d r a t s   f � r e   d e t   d a t u m e t 
 E x e m p e l :   * . z i p > 1 G ;   < 2 0 1 2 - 0 1 - 2 1  S e   h j � l p   f � r   f l e r   a l t e r n a t i v .  U T F - 8 � * * F � l j a n d e   a n v � n d a r s t a t i s t i k s d a t a   s k i c k a s   a n o n y m t   t i l l   W i n S C P . * * 
 
 U n d e r   t i d e n   k a n   a n n a n   s t a t i s t i k   s a m l a s   i n ,   k o m   g � r n a   t i l l b a k a   s e n a r e   f � r   a t t   k o n t r o l l e r a   e l l e r   k o n s u l t e r a   h j � l p e n . \ D e t   f i n n s   i n g e n   d a t a   i n s a m l a d   f � r   a n v � n d a r s t a t i s t i k   � n n u .   F � r s � k   i g e n   s e n a r e   e l l e r   s e   H j � l p .  � p p n a   w e b b p l a t s k a t a l o g   ' % s '  � p p n a r   a r b e t s y t a   ' % s '  S e n a s t e   a r b e t s y t o r  M i n   a r b e t s y t a - A r b e t s y t a   ' % s '   k o m m e r   a t t   s p a r a s   a u t o m a t i s k t .  A r b e t s y t a :   % s � * * � v e r f � r i n g s b e k r � f t e l s e   a v s t � n g d * * 
 
 D u   h a r   v a l t   a t t   i n t e   v i s a   d i a l o g r u t a n   f � r   � v e r f � r i n g s a l t e r n a t i v   n � s t a   g � n g .   K l i c k a   h � r   f � r   a t t   � n g r a .  F � r i n s t � l l n i n g a r 	 A v s l u t a d e u % s 
 
 D e t   u p p s t o d   n � g r a   f e l   v i d   k r y p t e r i n g e n   a v   l � s e n o r d   m e d   h j � l p   a v   e t t   n y t t   h u v u d l � s e n o r d   e l l e r   d e k r y p t e r a   l � s e n o r d . W i n S C P   � r   e n   p o p u l � r   g r a t i s   S F T P -   o c h   F T P - k l i e n t   f � r   W i n d o w s ,   e n   k r a f t f u l l   f i l h a n t e r a r e   s o m   k o m m e r   a t t   f � r b � t t r a   d i n   p r o d u k t i v i t e t .   D e n   s t � d e r   � v e n   l o k a l t   l � g e   o c h   F T P S - ,   S 3 - ,   S C P -   o c h   W e b D A V - p r o t o k o l l .   P o w e r - a n v � n d a r e   k a n   a u t o m a t i s e r a   W i n S C P   m e d   h j � l p   a v   . N E T - m o n t e r i n g . 	 L a d d a r . . . * % s 
 
 K l i c k a   h � r   f � r   a t t   s e   v a d   s o m   � r   n y t t . # % d   s l �   u p p   l � n k a r   o c h   l � s e r   k a t a l o g  K a n   i n t e   v i s a  A n v � n d n i n g : 5 N a m n   p �   w e b b p l a t s   e l l e r   d i r e k t   s e s s i o n s s p e c i f i k a t i o n . ; � p p n a   s e s s i o n   i   e t t   n y t t   f � n s t e r ,   � v e n   o m   % A P P %   k � r s   r e d a n . % � p p n a r   f j � r r f i l   i   d e n   i n t e r n a   e d i t o r . ) S y n k r o n i s e r a s   i n n e h � l l e t   i   t v �   k a t a l o g e r . - S t a r t a r   f u n k t i o n e n   h � l l   f j � r r k a t a l o g   a k t u e l l . / S t a r t a r   o p e r a t i o n   u t a n   a t t   v i s a   a l t e r n a t i v r u t a . @ K o n s o l   ( t e x t )   l � g e .   S t a n d a r d l � g e ,   n � r   d e n   a n r o p a s   m e d   % A P P % . c o m . b K � r   b a t c h s k r i p t f i l .   O m   s k r i p t e t   i n t e   s l u t a r   m e d   ' e x i t ' - k o m m a n d o t ,   n o r m a l t   i n t e r a k t i v t   l � g e   f � l j e r .  K � r   l i s t a   m e d   s k r i p t k o m m a n d o n . + S k i c k a r   l i s t a   m e d   p a r a m e t r a r   t i l l   s k r i p t e t . # S � k v � g   t i l l   k o n f i g u r a t i o n s   I N I - f i l . D K o n f i g u r e r a r   i n s t � l l n i n g a r   m e d   h j � l p   a v   R A W - f o r m a t   s o m   i   e n   I N I - f i l . f U p p d a t e r i n g s i n s t � l l n i n g a r   a v   w e b b p l a t s e r   s o m   m a t c h a r   e n   m a s k   m e d   h j � l p   a v   r a w - f o r m a t   s o m   i   e n   I N I - f i l . # A k t i v e r a r   s e s s i o n l o g g n i n g   t i l l   f i l . E L o g g i n g s n i v �   ( 0 . . 2 ) ,   l � g g a   t i l l   *   f � r   a t t   a k t i v e r a   l � s e n o r d s l o g g n i n g .   A k t i v e r a r   X M L - l o g g n i n g   t i l l   f i l . 8 G r u p p e r a   a l l a   X M L - l o g e l e m e n t   s o m   t i l l h � r   s a m m a   k o m m a n d o .  S S H   p r i v a t   n y c k e l f i l ) F i n g e r a v t r y c k   a v   s e r v e r n s   S S H - v � r d n y c k e l .  T L S / S S L - k l i e n t c e r t i f i k a t f i l .  P a s s i v t   l � g e   ( F T P - p r o t o k o l l ) . ! I m p l i c i t   T L S / S S L   ( F T P - p r o t o k o l l ) . ! E x p l i c i t   T L S / S S L   ( F T P - p r o t o k o l l ) .  S e r v e r n   s v a r a d e   m e d   t i m e o u t . Q K o n f i g u r e r a r   a l l a   s e s s i o n s i n s t � l l n i n g a r   m e d   h j � l p   a v   R A W - f o r m a t   s o m   i   e n   I N I   f i l . + H e m s i d a   f � r   f � r f r � g n i n g a r   o m   u p p d a t e r i n g a r .  S k r i v e r   u t   d e n n a   a n v � n d n i n g . � K o n v e r t e r a r   p r i v a t   n y c k e l   t i l l   . p p k - f o r m a t   e l l e r   r e d i g e r a r   n y c k e l .   A n v � n d   % s   f � r   a t t   a n g e   u t d a t a f i l .   A n v � n d   % s   f � r   a t t   � n d r a   e l l e r   s t � l l a   i n   l � s e n o r d s f r a s .   A n v � n d   % s   f � r   a t t   � n d r a   e l l e r   s t � l l a   i n   k o m m e n t a r .   A n v � n d   % s   f � r   a t t   l � g g a   t i l l   c e r t i f i k a t . $ A n g e   l � s e n f r a s   f � r   a t t   s p a r a   n y c k e l : ) M a t a   � t e r   i n   l � s e n o r d s f r a s   f � r   v e r i f i e r a :  N y c k e l   s p a r a d   t i l l   " % s " . D F i n g e r a v t r y c k   f � r   s e r v e r   T L S / S S L - c e r t i f i k a t   ( e n d a s t   F T P S - p r o t o k o l l ) .  G e r   e t t   n a m n   t i l l   s e s s i o n e n � U p p d a t e r a r   f j � r r p a n e l e n   f � r   a l l a   i n s t a n s e r   a v   W i n S C P .   O m   e n   s e s s i o n   ( o c h   e v e n t u e l l t   e n   s � k v � g )   a n g e s ,   u p p d a t e r a r   e n d a s t   i n s t a n s e n   m e d   d e n   s e s s i o n e n   ( o c h   s � k v � g e n ) . ? A k t i v e r a r   l o g g r o t a t i o n   o c h   e v e n t u e l l t   r a d e r i n g   a v   g a m l a   l o g g a r .  L � s e n o r d e t   h a r   � n d r a t s .  � p p n a   & m � l m a p p e n  � p p n a   & n e d l a d d a d   f i l � * * K r y p t e r i n g s n y c k e l   g e n e r e r a d e s . * * 
 
 D u   b � r   s � k e r h e t s k o p i e r a   d e n   g e n e r e r a d e   k r y p t e r i n g s n y c k e l n .   O m   d u   f � r l o r a r   d e n   k a n   d u   i n t e   l � s a   d i n a   k r y p t e r a d e   f i l e r . > � p p n a   p l a t s p r o f i l   " % s " . | L o k a l   k a t a l o g : 
     % s | F j � r r k a t a l o g : 
     % s : S k r i v e r   u t   e n   l i s t a   � v e r   c h i f f e r   o c h   a l g o r i t m e r   s o m   s t � d s . H K o n f i g u r e r a r   � v e r f � r i n g s i n s t � l l n i n g a r   m e d   e t t   r � f o r m a t   s o m   i   e n   I N I - f i l . D ! E   e x p a n d e r a r   t i l l   s e r i a l i s e r a d e   a n s l u t n i n g s d a t a   f � r   a k t u e l l   s e s s i o n   F E t t   l � s e n o r d   f � r   e n   k r y p t e r a d   p r i v a t   n y c k e l   e l l e r   e t t   k l i e n t c e r t i f i k a t B T r y c k   p �   ' N e j '   f � r   a t t   a k t i v e r a   a u t o m a t i s k   s p a r n i n g   a v   a r b e t s y t a n . ( V � l j e r   d e n   a n g i v n a   f i l e n   i   f i l p a n e l e r n a . � * * R e d i g e r a   t e r m i n a l i n s t � l l n i n g a r   i   P u T T Y . * * 
 
 P u T T Y   k o m m e r   a t t   s t a r t a s .   R e d i g e r a   t e r m i n a l i n s t � l l n i n g a r   f � r   e n   t i l l f � l l i g   w e b b p l a t s   % s .   W i n S C P   k o m m e r   i h � g   d e s s a   i n s t � l l n i n g a r   e f t e r   a t t   d u   s t � n g e r   P u T T Y .  T e r m i n a l i n s t � l l n i n g a r   f � r   % s 8 E t t   a l t e r n a t i v t   s � t t   a t t   t i l l h a n d a h � l l a   e t t   a n v � n d a r n a m n 4 E t t   a l t e r n a t i v t   s � t t   a t t   t i l l h a n d a h � l l a   e t t   l � s e n o r d ! A l l a   p r o m p t e r   a v b r y t s   a u t o m a t i s k t R T i l l � t e r   s t r e a m i n g   a v   f i l e r   t i l l   s t d o u t   ( o c h   o m d i r i g e r a r   s t a t u s u t d a t a   t i l l   s t d e r r ) & T i l l � t e r   s t r � m n i n g   a v   f i l e r   f r � n   s t d i n  T a r   b o r t . . .  T a c k   f � r   a t t   d u   k � p t e   W i n S C P . 2 L � s   m e r   o m   a t t   g �   � v e r   f r � n   k l a s s i s k   i n s t a l l a t i o n .  I g n o r e r a  L � s   a l l a   l � s e n o r d   f r � n   f i l e r  D i n   v e r s i o n :   % s  W I N _ F O R M S _ S T R I N G S          % s   f i l   ' % s '   t i l l   % s :  % s   % d   f i l e r   t i l l   % s :      l o k a l   k a t a l o g  f j � r r k a t a l o g    F l y t t a 	 s l � p p   m � l            T a r   b o r t  S t � l l e r   i n   i n s t � l l n i n g a r  T e m p o r � r   k a t a l o g 
 N y   k a t a l o g     	 A v m a r k e r a  M a r k e r a  % d   f i l  % d   f i l e r 
 % d   k a t a l o g  % d   k a t a l o g e r  % d   s y m b o l i s k   l � n k  % d   s y m b o l i s k a   l � n k a r    % s   E g e n s k a p e r  % s ,   . . .   E g e n s k a p e r  A n g e   g i l t i g t   g r u p p n a m n .  A n g e   g i l t i g t   � g a r n a m n .  T i l l b a k a   t i l l   % s  F r a m � t   t i l l   % s      A n s l u t n i n g s t i d  K o m p r i m e r i n g   ( % s )      I n f o r m a t i o n   o m   v a l d   f i l     P � p p n a   s p a r a d   s e s s i o n   ' % s '   ( h � l l   n e r e   S H I F T   f � r   a t t   � p p n a   s e s s i o n   i   n y t t   f � n s t e r )    L i c e n s   f � r   % s                � p p n a   k a t a l o g  H a n t e r a   b o k m � r k e n             
 R a d :   % d / % d 
 K o l u m n :   % d  T e c k e n :   % d   ( 0 x % . 2 x )  � n d r a d  K a n   i n t e   h i t t a   s t r � n g e n   ' % s ' .  T o t a l t   a n t a l   e r s � t t n i n g a r :   % d  G �   t i l l   r a d 
 R a d n u m m e r :  O g i l t i g t   r a d n u m m e r .  R e d i g e r a   l � n k / g e n v � g  L � g g   t i l l   l � n k / g e n v � g  I n t e   a n s l u t e n  A n s l u t e r . . .  V � l j   f l i k e n   ' % s '  L � g g   t i l l   p l a t s p r o f i l  P l a t s p r o f i l n a m n :    F l y t t a   p l a t s p r o f i l  N y t t   k a t a l o g n a m n :  S p a r a   s e s s i o n   s o m  & S p a r a   s e s s i o n   s o m : $ S p a r a   & l � s e n o r d   ( r e k o m m e n d e r a s   i n t e )    K � r   e g e t   k o m m a n d o               5 % s ,   % d   p t 
 T h e   Q u i c k   B r o w n   F o x   J u m p s   O v e r   T h e   L a z y   D o g  O k � n d  B e r � k n a   k a t a l o g s t o r l e k        A l l m � n n a   i n s t � l l n i n g a r  L a g r a d e   s e s s i o n e r 
 C a c h e m i n n e  K o n f i g u r a t i o n e n s   I N I - f i l  S l u m p t a l s f r �   f i l  V � l j   l o k a l   k a t a l o g .  F l y t t a r      F l y t t a  H � l l   f j � r r k a t a l o g e n   u p p d a t e r a d % B e h � l l e r   f j � r r k a t a l o g e n   u p p d a t e r a d . . .  T e m p o r � r a   k a t a l o g e r  N y   f i l  R e d i g e r a   f i l  & S k r i v   f i l n a m n : ( D u p l i c a t e   f i l e   ' % s '   t o   r e m o t e   d i r e c t o r y : ' D u p l i c a t e   % d   f i l e s   t o   r e m o t e   d i r e c t o r y :  D u b b l e r a  K o p i e r a r  L � g g   t i l l   e g e t   k o m m a n d o  R e d i g e r a   e g e t   k o m m a n d o  L  F          H � & m t a   f l e r . . .  V � l j   e d i t o r a p p l i k a t i o n . 0 K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s   i   % s   a v   % s , L � g g   t i l l   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g + R e d i g e r a   f � r i n s t � l l d   � v e r f � r i n g s i n s t � l l n i n g 	 S & t a n d a r d  & K o n f i g u r e r a . . .  E g & e t . . .  E g e t   k o m m a n d o  L � g g   t i l l   e d i t o r  R e d i g e r a   e d i t o r  % s ,   B a s e r a s   p �   % s   v e r s i o n   % s  & � p p n a    E n d a s t   & s a m m a   s t o r l e k   N u m b e r   o f   L i c e n s e s :   % s | U n l i m i t e d  P r o d u c t   I D :   % s  % s   ( E x p i r a t i o n   o n   % s )  % s       E d u c a t i o n a l   L i c e n s e  H � m t a r   e g e n s k a p e r    S S H   i m p l e m e n t a t i o n  K r y p t e r i n g s a l g o r i t m  K o m p r i m e r i n g  F i l � v e r f � r i n g s p r o t o k o l l  K a n   � n d r a   r � t t i g h e t e r  K a n   � n d r a   � g a r e / g r u p p  K a n   k � r a   g o d t y c k l i g t   k o m m a n d o " K a n   s k a p a   s y m b o l i s k   l � n k / h � r d   l � n k  K a n   s l �   u p p   a n v � n d a r g r u p p e r  K a n   d u b b l e r a   f j � r r f i l e r   $ � v e r f � r i n g s l � g e   f � r   r e n   t e x t   ( A S C I I ) $ K a n   k o n t r o l l e r a   t i l l g � n g l i g t   u t r y m m e  T o t a l t   a n t a l   b y t e s   p �   e n h e t  L e d i g t   a n t a l   b y t e s   p �   e n h e t   T o t a l t   a n t a l   b y t e s   f � r   a n v � n d a r e  L e d i g a   b y t e s   f � r   a n v � n d a r e  B y t e s   p e r   a l l o k e r i n g s e n h e t  O k � n d " H i t t a   P u T T Y / T e r m i n a l k l i e n t   k � r b a r a P P u T T Y / T e r m i n a l k l i e n t   k � r b a r a | % s | K � r b a r a   f i l e r   ( * . e x e ) | * . e x e | A l l a   f i l e r   ( * . * ) | * . *  % s   a v   % s | N / A  J � m f � r  S y n k r o n i s e r a r  A u t e n t i s e r i n g s b a n e r * I N I - f i l   ( * . i n i ) | * . i n i | A l l a   f i l e r   ( * . * ) | * . * ) V � l j   f i l   a t t   e x p o r t e r a   i n s t � l l n i n g a r   t i l l  S & e n a s t e :   % s  S & e n a s t e  B e r � k n a r   f i l k o n t r o l l s u m m a  K a n   b e r � k n a   f i l k o n t r o l l s u m m a  O k � n d  P r o t o k o l l   s o m   a n v � n d s    O s � k e r   a n s l u t n i n g  S � k e r   a n s l u t n i n g   ( % s )  E n d a s t   p r o t o k o l l k o m m a n d o n  F j � r r s y s t e m  K r y p t o g r a f i s k t   p r o t o k o l l      M i n a   d o k u m e n t 	 S k r i v b o r d    K o m m a n d o  S � t t   t i l l   s & t a n d a r d                            V � l j   l o k a l   p r o x y a p p l i k a t i o n � M � n s t e r : 
 \ n   f � r   n y   r a d 
 \ r   f � r   v a g n r e t u r 
 \ t   f � r   t a b b 
 \ x X X   f � r   h e x a d e c i m a l   a s c i i k o d 
 \ \   f � r   b a c k s l a s h 
 % v � r d   u t � k a s   t i l l   v � r d n a m n 
 % p o r t   u t � k a s   t i l l   p o r t n u m m e r 
 % u a n v � n d a r e   u t � k a s   t i l l   p r o x y a n v � n d a r n a m n 
 % l � s e n   u t � k a s   t i l l   p r o x y l � s e n o r d 
 % %   f � r   p r o c e n t t e c k e n = W e b b p l a t s k a t a l o g   e l l e r   a r b e t s y t a   m e d   n a m n e t   ' % s '   f i n n s   r e d a n . E � r   d u   s � k e r   a t t   d u   v i l l   r a d e r a   s e s s i o n s k a t a l o g   ' % s '   m e d   % d   s e s s i o n e r ? $ K a n   i n t e   r a d e r a   s p e c i a l s e s s i o n   ' % s ' .  S k a p a   s e s s i o n s k a t a l o g  N y t t   k a t a l o g n a m n :    H o w   t o   p u r c h a s e   a   l i c e n s e . . .  M � l f j � r r & s � k v � g : * * V i l l   d u   � p p n a   e n   s e p a r a t   s k a l s e s s i o n   f � r   a t t   d u p l i c e r a   % s ? * * 
   
 N u v a r a n d e   s e s s i o n   s t � d e r   i n t e   d i r e k t   d u p l i c e r i n g   a v   f j � r r s e s s i o n   % s .   E n   s e p a r a t   s k a l s e s s i o n   k a n   � p p n a s   f � r   a t t   b e a r b e t a   d u p l i c e r i n g e n .   A l t e r n a t i v t   k a n   d u   d u p l i c e r a   % s   v i a   l o k a l   t e m p o r � r   k o p i a .  f i l ( e r ) | k a t a l o g ( e r )  E d i t o r  % s   d o l d  % s   f i l t r e r a d  F i l t e r � A k t u e l l   s e s s i o n   t i l l � t e r   e n d a s t   f � r � n d r i n g   a v   U I D   � g a n d e t .   D e t   v a r   i n t e   m � j l i g t   a t t   l � s a   U I D   f r � n   k o n t o n a m n e t   " % s " .   S p e c i f i c e r a   U I D   e x p l i c i t   i s t � l l e t .    � v e r f � r   i   & b a k g r u n d e n  % s   ( l � g g   t i l l   i   � v e r f � r i n g s k � )  I n g e n  V � l j   k o r t k o m m a n d o  K o r & t k o m m a n d o : 
 O b e g r � n s a t  H u v u d l � s e n o r d  & N u v a r a n d e   h u v u d l � s e n o r d :  N & y t t   h u v u d l � s e n o r d :  U p p r e p a   h u v u d l � s e n o r d : - S p a r a   & l � s e n o r d   ( s k y d d a s   g e n o m   h u v u d l � s e n o r d ) 	 L e t a   i   % s  S � k 	 S � k e r   . . .  K l a r . 	 A v b r u t e n .    & S t a r t  & S t o p p  S p a r a   & l � s e n o r d  A v b r y t e r . . .  K o d n i n g :   % s c F i l e n   h a r   � n d r a t s .   � n d r i n g a r   k o m m e r   a t t   g �   f � r l o r a d e ,   o m   f i l e n   l a d d a s   m e d   a n n a n   k o d n i n g .   F o r t s � t t a ? F � r   d u   s � k e r   p �   a t t   d u   v i l l   t a   b o r t   a r b e t s y t a n   ' % s '   m e d   % d   s e s s i o n ( e r ) ?    S p a r a   a r b e t s y t a   s o m  & S p a r a   a r b e t s y t a   s o m : $ S p a r a   & l � s e n o r d   ( r e k o m m e n d e r a s   i n t e ) . S p a r a   & l � s e n o r d   ( s o m   s k y d d a s   a v   h u v u d l � s e n o r d )  S p a r a   & l � s e n o r d Q � p p n a   a r b e t s y t a   ' % s '   ( h � l l   n e r   S h i f t   f � r   a t t   � p p n a   a r b e t s y t a n   i   e t t   n y t t   f � n s t e r )  & � p p n a   k a t a l o g U � p p n a   w e b b p l a t s k a t a l o g   ' % s '   ( h � l l   n e r   S h i f t   f � r   a t t   � p p n a   k a t a l o g   i   e t t   n y t t   f � n s t e r )    & S k a p a   g e n v � g   p �   s k r i v b o r d e t , A k t i v e r a   & a u t o m a t i s k t   s p a r a n d e   a v   a r b e t s y t a n  H � m t a  � v e r f � r  H � m t a  � v e r f � r ) % s   f i l   ' % s '   t i l l   % s   o c h   t a   b o r t   o r i g i n a l : + % s   % d   f i l e r   t i l l   % s   o c h   t a   b o r t   o r i g i n a l e n :  H � m t a   o c h   t a   b o r t  � v e r f � r   o c h   t a   b o r t  K �  I m p o r t e r a   w e b b p l a t s e r - F e l   v i d   l a d d n i n g   a v   f i l   ' % s '   m e d   ' % s '   k o d n i n g                        F e l   v i d   l a d d n i n g   a v   f i l   ' % s ' .  � t e r g � r   t i l l   ' % s '   k o d n i n g . ) V � l j   f i l   a t t   i m p o r t e r a   k o n f i g u r a t i o n   f r � n  S � k :   % s  ( t r y c k   p �   t a b b   f � r   n � s t a )  � v e r f � r  H � m t a r  % d   i   k � �M � n s t e r : 
 ! !   e x p a n d e r a r   t i l l   u t r o p s t e c k e n 
 ! /   e x p a n d e r a r   t i l l   a k t u e l l   f j � r r s � k v � g 
 ! @   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   v � r d n a m n 
 ! U   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   a n v � n d a r n a m n 
 ! P   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   l � s e n o r d 
 ! #   e x p a n d e r a r   t i l l   a k t u e l l   s e s s i o n s   p o r t n u m m e r 
 ! N   e x p a n d e r a r   t i l l   a k t u e l l t   s e s s i o n s n a m n 
 ! ? p r o m p t [ \ ] ? d e f a u l t !   e x p a n d e r a r   t i l l   a n v � n d a r v a l t   v � r d e   m e d   g i v e n   p r o m p t   o c h   s t a n d a r d   ( a l t e r n a t i v t   \   u n d v i k e r   e s c a p e ) 
 ! ` c o m m a n d `   e x p a n d e r a r   t i l l   u t d a t a   a v   l o k a l t   k o m m a n d o  N y   w e b b p l a t s  K a t a l o g   w e b b p l a t s 	 A r b e t s y t a 8 D u   r e d i g e r a r   e n   w e b b p l a t s .   V i l l   d u   s p a r a   d i n a   � n d r i n g a r ? 	 & K a t a l o g :  < i n g e n >  S k a l  S C P / S k a l  E d i t o r   2 � t e r s t � l l   s e s s i o n   ( p a n e l )   f � r g   t i l l   s y s t e m s t a n d a r d  F & l e r   f � r g e r . . .  V � l j   f � r g   p �   s e s s i o n   ( p a n e l )  A & v l � g s n a   B O M   o c h   E O F   t e c k e n  A & v l � g s n a   B O M   t e c k e n T L i c e n s a v t a l e n   f � r   f � l j a n d e   p r o g r a m   ( b i b l i o t e k )   � r   d e l   a v   a p p l i k a t i o n e n s   l i c e n s a v t a l .  V i s a   l i c e n s  T o o l b a r 2 0 0 0   l i b r a r y   % s  C o p y r i g h t   �   J o r d a n   R u s s e l l ! h t t p s : / / j r s o f t w a r e . o r g / t b 2 k d l . p h p  T B X   l i b r a r y   % s , C o p y r i g h t   �   A l e x   A .   D e n i s o v   a n d   c o n t r i b u t o r s ! h t t p s : / / g i t h u b . c o m / p l a s h e n k o v / T B X ' F i l e m a n a g e r   T o o l s e t   l i b r a r y   V e r s i o n   2 . 6  C o p y r i g h t   �   I n g o   E c k e l  J E D I   C o d e   L i b r a r y   ( J C L )   % s  h t t p s : / / j c l . d e l p h i - j e d i . o r g /  P n g C o m p o n e n t s   1 . 9 & C o p y r i g h t   �   U w e   R a a b e   a n d   M a r t i j n   S a l y ) h t t p s : / / g i t h u b . c o m / U w e R a a b e / P n g C o m p o n e n t s 	 S p a r a r . . .    S v e n s k   � v e r s � t t n i n g :  C o p y r i g h t   % s  F i l :  S � k v � g :  L � s n i n g 
 U p p l � s n i n g 	 & S t a n d a r d % � t e r s t � l l   e d i t o r n s   f � r g   t i l l   s t a n d a r d  V � l j   n � g o n   f � r g   t i l l   e d i t o r n  S p a r a   k o n v e r t e r a d   p r i v a t   n y c k e l ; P u T T Y   p r i v a t   n y c k e l f i l e r   ( * . p p k ) | * . p p k | A l l a   f i l e r   ( * . * ) | * . * / P r i v a t   n y c k e l   k o n v e r t e r a d   o c h   s p a r a d   t i l l   ' % s ' .    S k a p a   f i l - U R L  S k a p a   s e s s i o n - U R L / k o d  U R L  S k r i p t  k o d  D i t t   k o m m a n d o   % d  T i p s   % d   a v   % d  T i p s % K � r   a n p a s s a d e   k o m m a n d o t   ' % s '   s o m   ' % s '  K o m m a n d o r a d s a r g u m e n t  K o m m a n d o r a d s a r g u m e n t   f � r   % s K E n   s e r v e r v � r d s n y c k e l   � r   o k � n d .   A n s l u t   m i n s t   e n   g � n g ,   i n n a n   d u   s k a p a r   k o d e n .  C : \ s k r i v b a r \ s � k v � g \ t i l l \ l o g g \  S k a p a   & k o d . . .  S k a p a   � v e r f � r i n g s k o d   " K � r   s k r i p t e t   m e d   e t t   k o m m a n d o   s o m :   C : \ s � k v � g \ t i l l \ s c r i p t \ s c r i p t . t x t  D i n   k o d   ! K o n f i g u r e r a   � v e r f � r i n g s a l t e r n a t i v  � v e r f � r   f i l e r c E t t   t e s t f i l l i s t a   a n v � n d s   e n d a s t ,   � v e r v � g   a t t   a n v � n d a   e n   f i l m a s k   f � r   a t t   v � l j a   f i l e r   f � r   � v e r f � r i n g .  S � k   e f t e r   u p p d a t e r i n g a r  L � g g   t i l l   u t � k n i n g $ A n g e   U R L   e l l e r   s � k v � g   t i l l   u t � k n i n g :     
 B l � d d r a . . . 	 V � l j   ' % s '  & P a u s a   i   s l u t e t  & S e s s i o n s l o g g f i l  V � l j   f i l   f � r   s e s s i o n s l o g g . 4 S e s s i o n s l o g g f i l a r   ( * . l o g ) | * . l o g | A l l a   f i l e r   ( * . * ) | * . *  A n v � n d a r s t a t i s t i k    & F i l t e r :  & K o p i e r a   t i l l   u r k l i p p  V � r d :   % s 
 V � r d n y c k e l :   % s  K & o p i e r a  & M a r k e r a   a l l t  K o r & t k o m m a n d o :                    A l l m � n t  A n s l u t e n 0 A n s l u t e n   m e d   % s .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .   * A n s l u t e n   m e d   % s ,   f � r m e d l a r   S S L - k o p p l i n g . . .  A n s l u t e r   t i l l   % s   . . .  L i s t n i n g   a v   k a t a l o g e r   l y c k a d  K o p p l a r   i f r � n   s e r v e r    s t a r t a r   n e r l a d d n i n g   a v   % s  N e r l a d d n i n g   l y c k a d   * F � r s � k e r   a t t   a n s l u t a   % s   g e n o m   F T P   p r o x y . . .                 � t e r f � r   l i s t n i n g   a v   k a t a l o g e r . . . 7 S S L - k o p p l i n g   u p p r � t t a d .   V � n t a r   p �   v � l k o m s t m e d d e l a n d e . . .  S S L - k o p p l i n g   u p p r � t t a d  S t a r t a r   � v e r f � r i n g   a v   % s  � v e r f � r i n g   l y c k a d     # H � m t a r   f i l i n f o r m a t i o n   f r a m g � n g s r i k t  H � m t a r   f i l i n f o r m a t i o n . . .  K u n d e   i n t e   h � m t a   f i l i n f o r m a t i o n                   5 K u n d e   i n t e   s k a p a   s o c k e t   i   d e n   a n g i v n a   p o r t i n t e r v a l l e t    K a n   i n t e   u p p r � t t a   S S L - k o p p l i n g   ' K u n d e   i n t e   � t e r f �   l i s t n i n g   a v   k a t a l o g e r     # K a n   i n t e   i n i t i a l i s e r a   S S L - b i b l i o t e k         , � v e r f � r i n g s t u n n e l   k a n   i n t e   � p p n a s .   O r s a k :   % s    K a n   i n t e   t o l k a   v � r d n a m n   " % s " > � t e r u p p t a g n i n g s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   s k r i v a   � v e r   f i l . I P a u s k o m m a n d o   s t � d s   i n t e   a v   s e r v e r ,   m e n   l o k a l   o c h   f j � r r f i l s t o r l e k   � r   l i k a . , O f � r m � g e n   a t t   s k i c k a   k o m m a n d o .   K o p p l a   i f r � n .    P e e r   c e r t i f i k a t   f � r k a s t a s    N e r l a d d n i n g   a v b r u t e n                      F i l e n   f i n n s   r e d a n          P r o x y   k r � v e r   a u t e n t i s e r i n g P N � d v � n d i g   a u t e n t i s e r i n g s t y p   r a p p o r t e r a d   a v   p r o x y s e r v e r   � r   o k � n d   e l l e r   s t � d s   i n t e % K a n   i n t e   a v g � r a   v � r d   t i l l   p r o x y s e r v e r ! K a n   i n t e   a n s l u t a   t i l l   p r o x y s e r v e r C B e g � r a n   f r � n   p r o x y   m i s s l y c k a d e s ,   k a n   i n t e   a n s l u t a   g e n o m   p r o x y s e r v e r                        T i m e o u t   d e t e k t e r a d .  � v e r f � r i n g   a v b r u t e n            K u n d e   i n t e   s � t t a   f i l p e k a r e  O k � n t   f e l   i   S S L - l a g r e t % K u n d e   i n t e   v e r i f i e r a   S S L - c e r t i f i k a t e t                                                            1 0 0     5 A n s l u t n i n g   m e d   p r o x y   e t a b l e r a d ,   u t f � r   h a n d s k a k n i n g . . .  k o n t r o l l a n s l u t n i n g  d a t a a n s l u t n i n g                            W I N _ V A R I A B L E $ C o p y r i g h t   �   2 0 0 0  2 0 2 5   M a r t i n   P r i k r y l  h t t p s : / / w i n s c p . n e t / # h t t p s : / / w i n s c p . n e t / e n g / d o c s / h i s t o r y    h t t p s : / / w i n s c p . n e t / f o r u m /  h t t p s : / / w i n s c p . n e t / u p d a t e s . p h p # h t t p s : / / w i n s c p . n e t / e n g / d o w n l o a d . p h p ! h t t p s : / / w i n s c p . n e t / e n g / d o n a t e . p h p + h t t p s : / / w i n s c p . n e t / e n g / d o c s / ? v e r = % s & l a n g = % s - h t t p s : / / w i n s c p . n e t / e n g / d o c s / % s ? v e r = % s & l a n g = % s ' h t t p s : / / w i n s c p . n e t / e n g / t r a n s l a t i o n s . p h p : h t t p s : / / w i n s c p . n e t / e n g / d o c s / s e a r c h . p h p ? v e r = % s & l a n g = % s & q = % s K h t t p s : / / w i n s c p . n e t / f o r u m / p o s t i n g . p h p ? m o d e = n e w t o p i c & v e r = % s & l a n g = % s & r e p o r t = % s " h t t p s : / / w i n s c p . n e t / e n g / u p g r a d e . p h p 8 h t t p s : / / w w w . m i c r o s o f t . c o m / s t o r e / a p p s / 9 p 0 p q 8 b 6 5 n 8 x ? c i d = % s   + h t t p s : / / w i n s c p . n e t / e n g / d o c s / m i c r o s o f t _ s t o r e 1 h t t p s : / / w i n s c p . n e t / u p d a t e n e w s . p h p ? s t o r e _ g e t _ i m g = 1                                             5 G e n e r a t e H t t p U r l . G e n e r a t e   & H T T P   U R L = G e n e r e r a   & H T T P - U R L ^ G e n e r a t e H t t p U r l . G e n e r a t e s   H T T P   U R L   o f   t h e   s e l e c t e d   f i l e = G e n e r e r a r   H T T P - U R L   f � r   d e n   v a l d a   f i l e n  G e n e r a t e H t t p U r l . U R L = U R L T G e n e r a t e H t t p U r l . T h e s e   o p t i o n s   a r e   s i t e - s p e c i f i c . = D e s s a   a l t e r n a t i v   � r   p l a t s s p e c i f i k a . 8 G e n e r a t e H t t p U r l . & W e b   r o o t   p a t h : = & W e b b s e r v e r n s   r o t s � k v � g : ( G e n e r a t e H t t p U r l . U s e   H T T P & S = A n v � n d   H T T P & S C G e n e r a t e H t t p U r l . & U R L   r o o t   p a t h   ( o p t i o n a l ) : = & U R L   r o t s � k v � g   ( v a l f r i ) : c G e n e r a t e H t t p U r l . & W e b   s e r v e r   h o s t n a m e   o v e r r i d e   ( o p t i o n a l ) : = � s i d o s � t t   w e b b s e r v e r n s   v � r d n a m n   ( v a l f r i ) : " G e n e r a t e H t t p U r l . O p t i o n s = A l t e r n a t i v $ G e n e r a t e H t t p U r l . D i s p l a y   U R L = V i s a   U R L > G e n e r a t e H t t p U r l . C o p y   U R L   t o   c l i p b o a r d = K o p i e r a   U R L   t i l l   u r k l i p p ? G e n e r a t e H t t p U r l . O p e n   U R L   i n   w e b   b r o w s e r = � p p n a   U R L   i   w e b b l � s a r e n ) C o m p a r e F i l e s . & C o m p a r e   F i l e s = & J � m f � r   f i l e r � C o m p a r e F i l e s . C o m p a r e s   t h e   s e l e c t e d   l o c a l   a n d   r e m o t e   p a t h   u s i n g   a n   e x t e r n a l   f i l e   c o m p a r i s o n   t o o l = J � m f � r   v a l d   l o k a l   o c h   f j � r r s � k v � g   m e d   h j � l p   a v   e t t   e x t e r n t   v e r k t y g   f � r   j � m f � r e l s e   a v   f i l e r  C o m p a r e F i l e s . O p t i o n s = A l t e r n a t i v C C o m p a r e F i l e s . S e l e c t   & f i l e   c o m p a r i s o n   t o o l : = V � l j   & j � m f � r e l s e v e r k t y g : ! C o m p a r e F i l e s . A u t o m a t i c = A u t o m a t i s k < V e r i f y F i l e C h e c k s u m . V e r i f y   & C h e c k s u m = V e r i f i e r a   & k o n t r o l l s u m m a � V e r i f y F i l e C h e c k s u m . C o m p a r e s   c h e c k s u m s   o f   t h e   s e l e c t e d   l o c a l   a n d   r e m o t e   f i l e = J � m f � r   k o n t r o l l s u m m o r   f � r   d e n   v a l d a   l o k a l a   o c h   f j � r r f i l e n 1 S e a r c h T e x t . & S e a r c h   f o r   T e x t . . . = & S � k   e f t e r   t e x t . . . � S e a r c h T e x t . S e a r c h e s   r e c u r s i v e l y   f o r   a   t e x t   i n   t h e   c u r r e n t   r e m o t e   d i r e c t o r y = S � k e r   r e k u r s i v t   e f t e r   e n   t e x t   i   d e n   a k t u e l l a   f j � r r k a t a l o g e n  S e a r c h T e x t . T e x t : = T e x t :  S e a r c h T e x t . F i l e   m a s k : = F i l m a s k : 2 Z i p U p l o a d . & Z I P   a n d   U p l o a d . . . = & Z I P   o c h   l a d d a   u p p . . .   � Z i p U p l o a d . P a c k s   t h e   s e l e c t e d   f i l e s   t o   a   Z I P   a r c h i v e   a n d   u p l o a d s   i t = P a k e t e r a r   d e   v a l d a   f i l e r n a   t i l l   e t t   Z I P - a r k i v   o c h   l a d d a r   u p p   d e t   $ Z i p U p l o a d . & A r c h i v e   n a m e : = & A r k i v n a m n : " Z i p U p l o a d . U s e   & 7 - z i p = A n v � n d   & 7 - z i p < Z i p U p l o a d . A r c h i v e   & t y p e   ( w i t h   7 - z i p ) : = A r k i v & t y p   ( m e d   7 - z i p ) : F Z i p U p l o a d . 7 - z i p   & p a t h   ( 7 z . e x e / 7 z a . e x e ) : = 7 - z i p   s � k v � g   ( 7 z . e x e / 7 z a . e x e ) :  Z i p U p l o a d . L o g g i n g = L o g g n i n g W K e e p L o c a l U p T o D a t e . & K e e p   L o c a l   D i r e c t o r y   u p   t o   D a t e . . . = & H � l l   l o k a l   k a t a l o g   u p p d a t e r a d . . . � K e e p L o c a l U p T o D a t e . P e r i o d i c a l l y   s c a n s   f o r   c h a n g e s   i n   a   r e m o t e   d i r e c t o r y   a n d   r e f l e c t s   t h e m   o n   a   l o c a l   d i r e c t o r y = S k a n n a r   p e r i o d i s k t   e f t e r   f � r � n d r i n g a r   i   e n   f j � r r k a t a l o g   o c h   � t e r s p e g l a r   d e m   p �   e n   l o k a l   k a t a l o g ' K e e p L o c a l U p T o D a t e . D i r e c t o r i e s = K a t a l o g e r h K e e p L o c a l U p T o D a t e . & W a t c h   f o r   c h a n g e s   i n   t h e   r e m o t e   d i r e c t o r y : = & T i t t a   e f t e r   f � r � n d r i n g a r   i   f j � r r k a t a l o g e n � K e e p L o c a l U p T o D a t e . . . .   & a n d   a u t o m a t i c a l l y   r e f l e c t   t h e m   o n   t h e   l o c a l   d i r e c t o r y : = . . .   & o c h   r e f l e k t e r a   d e m   a u t o m a t i s k t   p �   d e n   l o k a l a   k a t a l o g e n : $ K e e p L o c a l U p T o D a t e . O p t i o n s = A l t e r n a t i v . K e e p L o c a l U p T o D a t e . & D e l e t e   f i l e s = & T a   b o r t   f i l e r < K e e p L o c a l U p T o D a t e . & B e e p   o n   c h a n g e = & S y s t e m l j u d   v i d   f � r � n d r i n g 6 K e e p L o c a l U p T o D a t e . C o n t i n u e   o n   & e r r o r = F o r t s � t t   v i d   & f e l A K e e p L o c a l U p T o D a t e . & I n t e r v a l   ( i n   s e c o n d s ) : = I n t e r v a l l   ( i   s e k u n d e r ) : & K e e p L o c a l U p T o D a t e . F i l e   & m a s k : = F i l m a s & k " K e e p L o c a l U p T o D a t e . L o g g i n g = L o g g n i n g 0 B a t c h R e n a m e . B a t c h   & R e n a m e . . . = B a t c h ,   & b y t   n a m n . . . w B a t c h R e n a m e . R e n a m e s   r e m o t e   f i l e s   u s i n g   a   r e g u l a r   e x p r e s s i o n = B y t e r   n a m n   p �   f j � r r f i l e r   m e d   h j � l p   a v   e t t   r e g u l j � r t   u t t r y c k  B a t c h R e n a m e . R e n a m e = B y t   n a m n j B a t c h R e n a m e . R e p l a c e   f i l e   n a m e   p a r t   m a t c h i n g   t h i s   p a t t e r n : = E r s � t t   d e l   a v   f i l n a m n   s o m   m a t c h a r   d e t t a   m � n s t e r :  B a t c h R e n a m e . w i t h : = m e d :  B a t c h R e n a m e . O p t i o n s = A l t e r n a t i v 4 B a t c h R e n a m e . & P r e v i e w   c h a n g e s = F � & r h a n d s v i s a   � n d r i n g a r  B a t c h R e n a m e . L o g g i n g = L o g g n i n g ? A r c h i v e D o w n l o a d . & A r c h i v e   a n d   D o w n l o a d . . . = & A r k i v e r a   o c h   h � m t a . . . A r c h i v e D o w n l o a d . P a c k s   t h e   s e l e c t e d   f i l e s   t o   a n   a r c h i v e ,   d o w n l o a d s   i t ,   a n d   o p t i o n a l l y   e x t r a c t s   t h e   a r c h i v e   t o   t h e   c u r r e n t   l o c a l   d i r e c t o r y = P a c k a r   d e   v a l d a   f i l e r n a   t i l l   e t t   a r k i v ,   l a d d a r   n e r   d e t   o c h   e x t r a h e r a r   e v e n t u e l l t   a r k i v e t   t i l l   d e n   a k t u e l l a   l o k a l a   k a t a l o g e n * A r c h i v e D o w n l o a d . & A r c h i v e   n a m e : = & A r k i v n a m n : ) A r c h i v e D o w n l o a d . A r c h i v e   & t y p e : = A r k i v & t y p :   A r c h i v e D o w n l o a d . P a c k i n g = P a c k n i n g A A r c h i v e D o w n l o a d . C u s t o m   a r c h i v e   & c o m m a n d : = A n p a s s a t   a r k i v & k o m m a n d o :   % A r c h i v e D o w n l o a d . E x t r a c t i n g = U p p a c k n i n g @ A r c h i v e D o w n l o a d . & E x t r a c t   a f t e r   d o w n l o a d = & P a c k   u p p   e f t e r   h � m t n i n g F A r c h i v e D o w n l o a d . U s e   & 7 - z i p   f o r   e x t r a c t i n g = A n v � n d   & 7 - z i p   f � r   u p p a c k n i n g L A r c h i v e D o w n l o a d . 7 - z i p   & p a t h   ( 7 z . e x e / 7 z a . e x e ) : = 7 - z i p   s � k v � g   ( 7 z . e x e / 7 z a . e x e ) :   A r c h i v e D o w n l o a d . L o g g i n g = L o g g n i n g m S y n c h r o n i z e A n o t h e r S e r v e r . & S y n c h r o n i z e   w i t h   A n o t h e r   R e m o t e   S e r v e r . . . = & S y n k r o n i s e r a   m e d   e n   a n n a n   f j � r r s e r v e r . . . S y n c h r o n i z e A n o t h e r S e r v e r . S y n c h r o n i z e s   a   d i r e c t o r y   o n   a n o t h e r   s e r v e r   ( o r   a n o t h e r   d i r e c t o r y   o n   t h i s   s e r v e r )   a g a i n s t   a   d i r e c t o r y   o n   t h i s   s e r v e r = S y n k r o n i s e r a r   e n   k a t a l o g   p �   e n   a n n a n   s e r v e r   ( e l l e r   e n   a n n a n   k a t a l o g   p �   d e n   h � r   s e r v e r n )   m o t   e n   k a t a l o g   p �   d e n   h � r   s e r v e r n j S y n c h r o n i z e A n o t h e r S e r v e r . S y n c h r o n i z e   d i r e c t o r y   f r o m   & t h i s   s e r v e r : = S y n k r o n i s e r a   k a t a l o g   f r � n   & d e n n a   s e r v e r : . S y n c h r o n i z e A n o t h e r S e r v e r . & D i r e c t o r y : = & K a t a l o g : K S y n c h r o n i z e A n o t h e r S e r v e r . . . .   t o   & a n o t h e r   s e r v e r : = . . .   t i l l   e n   & a n n a n   s e r v e r : , S y n c h r o n i z e A n o t h e r S e r v e r . & S e s s i o n : = & S e s s i o n : Y S y n c h r o n i z e A n o t h e r S e r v e r . & P r o m p t   f o r   s e s s i o n   p a s s w o r d = & F r � g a   e f t e r   l � s e n o r d   f � r   s e s s i o n e n . S y n c h r o n i z e A n o t h e r S e r v e r . D i & r e c t o r y : = K a & t a l o g : + S y n c h r o n i z e A n o t h e r S e r v e r . O p t i o n s = A l t e r n a t i v 5 S y n c h r o n i z e A n o t h e r S e r v e r . & D e l e t e   f i l e s = & T a   b o r t   f i l e r A S y n c h r o n i z e A n o t h e r S e r v e r . & P r e v i e w   c h a n g e s = F � & r h a n d s v i s a   � n d r i n g a r   = S y n c h r o n i z e A n o t h e r S e r v e r . C o n t i n u e   o n   & e r r o r = F o r t s � t t   v i d   & f e l ) S y n c h r o n i z e A n o t h e r S e r v e r . L o g g i n g = L o g g n i n g                             " S k a l t i l l � g g e t   � r   i n t e   i n s t a l l e r a t . 7 S k a l t i l l � g g e t   � r   i n s t a l l e r a t ,   m e n   d e t   h a r   i n t e   l a d d a t s . % S k a l t i l l � g g e t   i n s t a l l e r a s   o c h   l a d d a s . E * * P u b l i k   n y c k e l   f � r   a t t   k l i s t r a   i n   i   O p e n S S H   a u t h o r i z e d _ k e y s - f i l e n : * * � * * I n s t a l l e r a   d e n   p u b l i k a   n y c k e l n   t i l l   i c k e - O p e n S S H   s e r v e r ? * * 
 
 I n s t a l l e r i n g   a v   d e n   p u l i k a   n y c k e l n   s t � d s   e n d a s t   f � r   O p e n S S H   s e r v e r   ( a u t h o r i z e d _ k e y s - f i l ) . 
 
 D i n   s e r v e r   � r   % s . ! I n s t a l l e r a r   p u b l i k   n y c k e l   " % s " . . .     * V � l j   n y c k e l   f � r   a t t   i n s t a l l e r a   t i l l   s e r v e r � P u T T Y   p r i v a t a   n y c k e l f i l e r   ( * . p p k ) | * . p p k | A l l a   p r i v a t a   n y c k e l f i l e r   ( * . p p k ; * . p e m ; * . k e y ; i d _ * ) | * . p p k ; * . p e m ; * . k e y ; i d _ * | A l l a   f i l e r   ( * . * ) | * . *  C h e c k l i s t   f � r   s y n k r o n i s e r i n g  S k r i v s k y d d a d  B e r � k n a r  S p a r a   s o m   & f � r i n s t � l l n i n g . . .  B y t   n a m n   p �   f l i k e n  & N y t t   f l i k n a m n :  S y n k r o n i s e r i n g e n   s l u t f � r d e s . � U p p l a d d a d e   f i l e r :   % s   ( % s ) | N e d l a d d a d e   f i l e r :   % s   ( % s ) | L o k a l a   f i l e r   r a d e r a d e :   % s | E x t e r n a   f i l e r   r a d e r a d e :   % s | J � m f � r e l s e t i d :   % s | S y n k r o n i s e r i n g s t i d :   % s 1 S k a l t i l l � g g   k a n   i n t e   f u n g e r a   p �   d e t   h � r   s y s t e m e t .  F i l f � r g � F � r   a t t   a k t i v e r a   a u t o m a t i s k a   u p p d a t e r i n g a r ,   s n � l l a   < a   h r e f = " % D O N A T E _ U R L % " > d o n e r a   t i l l   W i n S C P - u t v e c k l i n g < / a >   e l l e r   % G E T _ I M G %   W i n S C P   f r � n   < a   h r e f = " % S T O R E _ U R L % " > M i c r o s o f t   S t o r e < / a > .  N y 	 S t a t i s t i k  R a w - w e b b p l a t s i n s t � l l n i n g a r  & L � g g   t i l l . . . " L � g g   t i l l   R a w - w e b b p l a t s i n s t � l l n i n g  & W e b b p l a t s i n s t � l l n i n g :  L a d d a   u p p   n y   l o k a l   f i l  L a d d a   n e r   n y   f j � r r f i l  L a d d a   u p p   u p p d a t e r a d   l o k a l   f i l  L a d d a   n e r   u p p d a t e r a d   f j � r r f i l  T a   b o r t   f � r � l d r a d   f j � r r f i l    T a   b o r t   f � r � l d r a d   l o k a l   f i l  K l i c k a   f � r   o m v � n t  & L o k a l  F & j � r r  & V � n s t e r  & H � g e r  K o p i e r a  F l y t t a  � p p n a  L o g g a   i n ] K l i c k a   f � r   a t t   � p p n a   e n   n y   l o k a l   f l i k . 
 H � l l   n e d   C t r l - t a n g e n t e n   f � r   a t t   � p p n a   e n   n y   f j � r r f l i k . x K l i c k a   f � r   a t t   � p p n a   n y   s e s s i o n   i   e n   n y   f j � r r f l i k . 
 H � l l   n e d   S k i f t - t a n g e n t e n   f � r   a t t   � p p n a   n y   s e s s i o n   i   e t t   n y t t   f � n s t e r . : % s 
 H � l l   n e d   C t r l - t a n g e n t e n   f � r   a t t   � p p n a   e n   n y   l o k a l   f l i k . q % d   n y c k e l f i l e r   i   % d   i m p o r t e r a d e   s e s s i o n e r   k o n v e r t e r a d e s   e l l e r   e r s a t t e s   m e d   b e f i n t l i g a   n y c k l a r   i   f o r m a t   s o m   s t � d s .  K a n   � n d r a   A C L  A C L :   
 & A n v � n d a r e  & A l l a  L � s   A C L 	 S k r i v   A C L  A l l m � n # B e h � v s   f � r   P o w e r S h e l l   7 . 3   o c h   n y a r e  - -   v a r n a   e f t e r   d e t t a   - -  3 D E S  B l o w f i s h  A E S  D E S  A r c f o u r  C h a C h a 2 0  A E S - G C M                    - -   v a r n a   e f t e r   d e t t a   - - ! D i f f i e - H e l l m a n   g r o u p   1   ( 1 0 2 4 - b i t ) " D i f f i e - H e l l m a n   g r o u p   1 4   ( 2 0 4 8 - b i t ) " D i f f i e - H e l l m a n   g r o u p   1 5   ( 3 0 7 2 - b i t ) " D i f f i e - H e l l m a n   g r o u p   1 6   ( 4 0 9 6 - b i t ) " D i f f i e - H e l l m a n   g r o u p   1 7   ( 6 1 4 4 - b i t ) " D i f f i e - H e l l m a n   g r o u p   1 8   ( 8 1 9 2 - b i t )  D i f f i e - H e l l m a n   g r u p p   u t b y t e  R S A - b a s e r a t   n y c k e l u t b y t e  E C D H   n y c k e l u t b y t e " N T R U   P r i m e   /   C u r v e 2 5 5 1 9   h y b r i d   k e x  M L - K E M   /   C u r v e 2 5 5 1 9   h y b r i d   k e x  M L - K E M   /   N I S T   E C D H   h y b r i d   k e x               � * * D e n n a   n y c k e l   i n n e h � l l e r   e t t   O p e n S S H - c e r t i f i k a t . * * 
 D e t   � r   i n t e   m e n i n g e n   a t t   d e n   s k a   l � g g a s   t i l l   i   f i l e n   O p e n S S H   a u t h o r i z e d _ k e y s . U M a t c h a n d e   c e r t i f i k a t   u p p t � c k t e s   i   ' % s '   o c h   l a d e s   t i l l   i   d e n   k o n v e r t e r a d e   n y c k e l f i l e n . ( R e d i g e r a   b e t r o d d   v � r d c e r t i f i k a t u t f � r d a r e ) L � g g   t i l l   b e t r o d d   v � r d c e r t i f i k a t u t f � r d a r e  & N a m n :  P u b l i k   & n y c k e l :   7 G i l t i g a   & v � r d a r   d e n n a   n y c k e l   � r   b e t r o d d   a t t   c e r t i f i e r a :  & B l � d d r a . . .   I n g e n   p u b l i k   n y c k e l   h a r   a n g e t t s . 2 V � l j   f i l   m e d   p u b l i k   n y c k e l   f � r   c e r t i f i k a t u t f � r d a r e 5 P u b l i c   n y c k e l f i l e r   ( * . p u b ) | * . p u b | A l l a   f i l e r   ( * . * ) | * . *                                           . D e t   g � r   i n t e   a t t   l a d d a   p u b l i k   n y c k e l   f r � n   ' % s ' # S i g n a t u r t y p e r   ( e n d a s t   R S A - n y c k l a r ) :  S H A - & 1 | S H A - & 2 5 6 | S H A - & 5 1 2 * I n g e t   v a l i d i t e t s u t t r y c k   h a r   k o n f i g u r e r a t s .  F e l   i   v a l i d i t e t s u t t r y c k . �* * S l u t a   v i s a   i n l o g g n i n g s d i a l o g r u t a n   a u t o m a t i s k t ? * *   B e k r � f t a   o m   d u   v e r k l i g e n   v i l l   a t t   W i n S C P   s l u t a r   v i s a   i n l o g g n i n g s d i a l o g r u t a n   a u t o m a t i s k t   v i d   s t a r t   o c h   n � r   d e n   s i s t a   s e s s i o n e n   s t � n g s . 
 
 O m   d u   � n d r a r   d i g   s e n a r e   k a n   d u   � t e r s t � l l a   d e t t a   i   I n s t � l l n i n g a r   p �   s i d a n   M i l j �   >   F � n s t e r . 
 
 F � r   a t t   � p p n a   i n l o g g n i n g s d i a l o g r u t a n   m a n u e l l t ,   g �   t i l l   F l i k a r   >   N y   f l i k   [ >   F j � r r f l i k ]   e l l e r   a n v � n d   m o t s v a r a n d e   k n a p p   i   v e r k t y g s f � l t e t . ' V � l j   f i l   a t t   i m p o r t e r a   w e b b p l a t s e r   f r � n    ( b � r j a   s k r i v a )  S � k  I n g a   s � k r e s u l t a t   h i t t a d e s .  R e d i g e r a   t a g g  L � g g   t i l l   t a g g  & N y c k e l :  & V � r d e   ( v a l f r i t t ) :                                   ? ! K   e x p a n d e r a r   t i l l   d e n   a k t u e l l a   s e s s i o n e n s   p r i v a t a   n y c k e l s � k v � g ' ! \   e x p a n d e r a r   t i l l   a k t u e l l   l o k a l   s � k v � g B I n s t a l l e r a r   d i n   p u b l i k a   n y c k e l   i   e n   s e r v e r s   a u k t o r i s e r a d e   n y c k l a r .                        a n   u n n a m e d   f i l e                       ' A n   u n s u p p o r t e d   o p e r a t i o n   w a s   a t t e m p t e d . $ A   r e q u i r e d   r e s o u r c e   w a s   u n a v a i l a b l e .  O u t   o f   m e m o r y .  A n   u n k n o w n   e r r o r   h a s   o c c u r r e d .                          N o   e r r o r   o c c u r r e d . - A n   u n k n o w n   e r r o r   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  % 1   w a s   n o t   f o u n d .  % 1   c o n t a i n s   a n   i n v a l i d   p a t h . = % 1   c o u l d   n o t   b e   o p e n e d   b e c a u s e   t h e r e   a r e   t o o   m a n y   o p e n   f i l e s .  A c c e s s   t o   % 1   w a s   d e n i e d . . A n   i n v a l i d   f i l e   h a n d l e   w a s   a s s o c i a t e d   w i t h   % 1 . < % 1   c o u l d   n o t   b e   r e m o v e d   b e c a u s e   i t   i s   t h e   c u r r e n t   d i r e c t o r y . 6 % 1   c o u l d   n o t   b e   c r e a t e d   b e c a u s e   t h e   d i r e c t o r y   i s   f u l l .  S e e k   f a i l e d   o n   % 1 5 A   h a r d w a r e   I / O   e r r o r   w a s   r e p o r t e d   w h i l e   a c c e s s i n g   % 1 . 0 A   s h a r i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 . 0 A   l o c k i n g   v i o l a t i o n   o c c u r r e d   w h i l e   a c c e s s i n g   % 1 .  D i s k   f u l l   w h i l e   a c c e s s i n g   % 1 . . A n   a t t e m p t   w a s   m a d e   t o   a c c e s s   % 1   p a s t   i t s   e n d .    I n v a l i d   h o u r   o f f s e t :   % d  I n v a l i d   d u r a t i o n   s t r i n g :   % s # H o u r   O f f s e t   p o r t i o n   o f   t i m e   i n v a l i d  I n v a l i d   d e c i m a l   s t r i n g :   ' ' % s ' ' 0 C a n n o t   c o n v e r t   s c i e n t i f i c   n o t a t i o n   t o   T B c d   v a l u e   C a n n o t   c o n v e r t   N A N   t o   T B c d   v a l u e ( I n v a l i d   B c d   P r e c i s i o n   ( % d )   o r   S c a l e   ( % d ) : C a n n o t   c o n v e r t   t o   T B c d :   s t r i n g   h a s   m o r e   t h a n   6 4   d i g i t s :   % s  % s   i s   n o t   a   v a l i d   h e x   s t r i n g  U n s u p p p o r t e d   v a r i a n t   t y p e   % d  v a r D i s p a t c h   t y p e   n o t   s u p p o r t e d  v a r E r r o r   t y p e   n o t   s u p p o r t e d  B C D   o v e r f l o w  % s   i s   n o t   a   v a l i d   B C D   v a l u e       ) % s   o n l y   s u p p o r t s   s i n k i n g   o f   m e t h o d   c a l l s ! & A t t e m p t i n g   t o   h o o k   c h i l d   w i n d o w s   t w i c e  S a v e   t h e   c u r r e n t   f i l e ? 0 O p e r a t i o n   n o t   s u p p o r t e d   b y   E d g e   W e b V i e w 2   c o n t r o l % F a i l e d   t o   c r e a t e   E d g e   b r o w s e r   c o n t r o l 2 T h e   u n d e r l y i n g   W e b V i e w 2   c o n t r o l   i s   n o t   i n i t i a l i z e d F I n t e r n a l   e r r o r :   d a t a   t y p e   k i n d   % s   c a n n o t   b e   c o n v e r t e d   t o   a n d   f r o m   t e x t + I n v o k a b l e   C l a s s   % s   i m p l e m e n t s   n o   i n t e r f a c e s  T y p e   c a n n o t   b e   c a s t   a s   V a r i a n t  I n t e r f a c e   % s   h a s   n o   R T T I 5 P a r a m e t e r   % s   o n   M e t h o d   % s   o f   I n t e r f a c e   % s   h a s   n o   R T T I  I n v a l i d   d a t e   s t r i n g :   % s  I n v a l i d   t i m e   s t r i n g :   % s  I n v a l i d   m i n u t e :   % d  I n v a l i d   m i l l i s e c o n d :   % d  I n v a l i d   f r a c t i o n a l   s e c o n d :   % f C 3 r d - l e v e l   c a c h e :   4   M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   8   M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e D 3 r d - l e v e l   c a c h e :   1 2   M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e D 3 r d - l e v e l   c a c h e :   1 8   M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e D 3 r d - l e v e l   c a c h e :   2 4   M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e  6 4 - B y t e   P r e f e t c h i n g  1 2 8 - B y t e   P r e f e t c h i n g e C P U I D   l e a f   2   d o e s   n o t   r e p o r t   c a c h e   d e s c r i p t o r   i n f o r m a t i o n ,   u s e   C P U I D   l e a f   4   t o   q u e r y   c a c h e   p a r a m e t e r s  I n v a l i d   M M F   n a m e   " % s " * T h e   M M F   n a m e d   " % s "   c a n n o t   b e   c r e a t e d   e m p t y  W i n 3 2   e r r o r :   % s   ( % u ) % s % s  L i b r a r y   n o t   f o u n d :   % s  F u n c t i o n   n o t   f o u n d :   % s . % s  N o   p a g e   l o a d e d  C a n n o t   r e g i s t e r   a   n i l   p r o v i d e r  I n v a l i d   s e r v i c e   p r o v i d e r   G U I D A I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   e n t r i e s ; D a t a   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   1 2 8   e n t r i e s < D a t a   T L B 1 :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   2 5 6   e n t r i e s ; D a t a   T L B 1 :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   e n t r i e s E D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   8   e n t r i e s C S h a r e d   2 n d - L e v e l   T L B :   4   K B y t e   p a g e s ,   4 - w a y   a s s o c i a t i v e ,   5 1 2   e n t r i e s D 3 r d - l e v e l   c a c h e :   5 1 2   K B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   1   M B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   2   M B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   1   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   2   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   4   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 3 r d - l e v e l   c a c h e :   1 . 5   M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   3   M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   6   M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   2   M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e   D 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e Z 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r Z 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r Z 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r X 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e s   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r C 2 n d - l e v e l   c a c h e :   2   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e A 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e A 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e ? 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e ? 2 n d - l e v e l   c a c h e :   2   M B y t e s ,   8 - w a y   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e D 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 2 n d - l e v e l   c a c h e :   1   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   1 2 8   e n t r i e s S I n s t r u c t i o n   T L B :   2   M B y t e   p a g e s ,   4 - w a y ,   8   e n t r i e s   o r   4   M B y t e   p a g e s ,   4 - w a y ,   4   e n t r i e s ; D a t a   T L B 0 :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   1 6   e n t r i e s 7 D a t a   T L B 0 :   4   K B y t e   p a g e s ,   4 - w a y   a s s o c i a t i v e ,   1 6   e n t r i e s 7 D a t a   T L B 0 :   4   K B y t e   p a g e s ,   f u l l y   a s s o c i a t i v e ,   1 6   e n t r i e s F D a t a   T L B 0 :   2   M B y t e   o r   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   e n t r i e s / D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   6 4   E n t r i e s 0 D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   1 2 8   E n t r i e s 0 D a t a   T L B :   4   K B y t e   a n d   4   M B y t e   p a g e s ,   2 5 6   E n t r i e s H 1 s t - l e v e l   d a t a   c a c h e :   1 6   K B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e H 1 s t - l e v e l   d a t a   c a c h e :   8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e I 1 s t - l e v e l   d a t a   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e I 1 s t - l e v e l   d a t a   c a c h e :   3 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e , T r a c e   c a c h e :   1 2   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e , T r a c e   c a c h e :   1 6   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e , T r a c e   c a c h e :   3 2   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e , T r a c e   c a c h e :   6 4   K - O p s ,   8 - w a y   s e t   a s s o c i a t i v e : I n s t r u c t i o n   T L B :   2 M / 4 M   p a g e s ,   f u l l y   a s s o c i a t i v e ,   8   e n t r i e s C 2 n d - l e v e l   c a c h e :   1   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e C 2 n d - l e v e l   c a c h e :   2   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   4   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   8   M B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   8   M B y t e ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e D 2 n d - l e v e l   c a c h e :   4   M B y t e s ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   6 M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 3 r d - l e v e l   c a c h e :   8 M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   1 2 M B y t e ,   1 2 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e C 3 r d - l e v e l   c a c h e :   1 6 M B y t e ,   1 6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e B 2 n d - l e v e l   c a c h e :   6 M B y t e ,   2 4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e * I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   3 2   E n t r i e s A I n s t r u c t i o n   T L B :   4   K B y t e   a n d   2   M B y t e   o r   4   M B y t e   p a g e s ,   6 4   E n t r i e s B I n s t r u c t i o n   T L B :   4   K B y t e   a n d   2   M B y t e   o r   4   M B y t e   p a g e s ,   1 2 8   E n t r i e s B I n s t r u c t i o n   T L B :   4   K B y t e   a n d   2   M B y t e   o r   4   M B y t e   p a g e s ,   2 5 6   E n t r i e s G I n s t r u c t i o n   T L B :   2 - M B y t e   o r   4 - M B y t e   p a g e s ,   f u l l y   a s s o c i a t i v e ,   7   e n t r i e s Y 3 r d   l e v e l   c a c h e :   5 1 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r W 3 r d   l e v e l   c a c h e :   1   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r W 3 r d   l e v e l   c a c h e :   2   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r W 3 r d   l e v e l   c a c h e :   4   M B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e ,   2   l i n e s   p e r   s e c t o r I 1 s t   l e v e l   d a t a   c a c h e :   3 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e P 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   3 2   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   1 9 2   K B y t e s ,   6 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   2 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   3 8 4   K B y t e s ,   6 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e U 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   s e c t o r e d   c a c h e ,   6 4 - b y t e   l i n e   s i z e X N o   2 n d - l e v e l   c a c h e   o r ,   i f   p r o c e s s o r   c o n t a i n s   a   v a l i d   2 n d - l e v e l   c a c h e ,   n o   3 r d - l e v e l   c a c h e E 2 n d - l e v e l   c a c h e :   1 2 8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   2 5 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e E 2 n d - l e v e l   c a c h e :   5 1 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e  F a i l e d   t o   o p e n   m u t e x  N u l l   d e s c r i p t o r A I n s t r u c t i o n   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   e n t r i e s @ I n s t r u c t i o n   T L B :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   2   e n t r i e s : D a t a   T L B :   4   K B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   e n t r i e s 9 D a t a   T L B :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   8   e n t r i e s ; D a t a   T L B 1 :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   e n t r i e s O 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   8   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e P 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e P 1 s t   l e v e l   i n s t r u c t i o n   c a c h e :   3 2   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e H 1 s t   l e v e l   d a t a   c a c h e :   8   K B y t e s ,   2 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e @ I n s t r u c t i o n   T L B :   4   M B y t e   p a g e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   4   e n t r i e s I 1 s t   l e v e l   d a t a   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   3 2   b y t e   l i n e   s i z e I 1 s t   l e v e l   d a t a   c a c h e :   1 6   K B y t e s ,   4 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e I 1 s t   l e v e l   d a t a   c a c h e :   2 4   K B y t e s ,   6 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e E 2 n d   l e v e l   c a c h e :   2 5 6   K B y t e s ,   8 - w a y   s e t   a s s o c i a t i v e ,   6 4   b y t e   l i n e   s i z e   
 E x e c u t a b l e  P a c k a g e  L i b r a r y 
 N e v e r B u i l d 
 D e s i g n O n l y  R u n O n l y  I g n o r e D u p U n i t s  D e l p h i   3   o r   C + +   B u i l d e r   3 	 U n d e f i n e d  C + +   B u i l d e r   4   o r   l a t e r  D e l p h i   4   o r   l a t e r  M a i n  W e a k  O r g W e a k  I m p l i c i t  F a i l e d   t o   c r e a t e   m u t e x    U n k n o w n  N a t i v e  G U I  C o n s o l e  O S / 2  P o s i x 
 R e s e r v e d   8  U N K N O W N  C O F F  C O D E V I E W  F P O  M I S C 	 E X C E P T I O N  F I X U P  O M A P _ T O _ S R C  O M A P _ F R O M _ S R C  A R M   L i t t l e - E n d i a n  T H U M B  A M 3 3  I B M   P o w e r P C   L i t t l e - E n d i a n  I B M   P o w e r P C   F P  I n t e l   6 4  M I P S 1 6  A L P H A 6 4  M I P S F P U 	 M I P S F P U 1 6  I n f i n e o n  C E F  E F I   B y t e   C o d e 
 A M D 6 4   ( K 8 )  M 3 2 R   l i t t l e - e n d i a n  C E E    P r o c e s s A f f i n i t y M a s k 
 C S D V e r s i o n  R e s e r v e d  E d i t L i s t  U n k n o w n 	 I n t e l   3 8 6  M I P S   l i t t l e - e n d i a n   R 3 0 0 0  M I P S   l i t t l e - e n d i a n   R 4 0 0 0  M I P S   l i t t l e - e n d i a n   R 1 0 0 0 0  M I P S   l i t t l e - e n d i a n   W C E   v 2 	 A l p h a _ A X P  S H 3   l i t t l e - e n d i a n  S H 3   D S P  S H 3 E   l i t t l e - e n d i a n  S H 4   l i t t l e - e n d i a n  S H 5  S i z e   o f   S t a c k   R e s e r v e  S i z e   o f   S t a c k   C o m m i t  S i z e   o f   H e a p   R e s e r v e  S i z e   o f   H e a p   C o m m i t  L o a d e r   F l a g s  N u m b e r   o f   R V A  V e r s i o n  G l o b a l F l a g s C l e a r  G l o b a l F l a g s S e t  C r i t i c a l S e c t i o n D e f a u l t T i m e o u t  D e C o m m i t F r e e B l o c k T h r e s h o l d  D e C o m m i t T o t a l F r e e T h r e s h o l d  L o c k P r e f i x T a b l e  M a x i m u m A l l o c a t i o n S i z e  V i r t u a l M e m o r y T h r e s h o l d  P r o c e s s H e a p F l a g s    S i z e   o f   U n i n i t i a l i z e d   D a t a  A d d r e s s   o f   E n t r y   P o i n t  B a s e   o f   C o d e  B a s e   o f   D a t a 
 I m a g e   B a s e  S e c t i o n   A l i g n m e n t  F i l e   A l i g n m e n t  O p e r a t i n g   S y s t e m   V e r s i o n  I m a g e   V e r s i o n  S u b s y s t e m   V e r s i o n  W i n 3 2   V e r s i o n  S i z e   o f   I m a g e  S i z e   o f   H e a d e r s  C h e c k S u m 	 S u b s y s t e m  D l l   C h a r a c t e r i s t i c s  I A T  D e l a y   l o a d   i m p o r t  C O M   r u n - t i m e  r e s e r v e d   [ % . 2 d ] 	 S i g n a t u r e  M a c h i n e  N u m b e r   o f   S e c t i o n s  T i m e   D a t e   S t a m p  S y m b o l s   P o i n t e r  N u m b e r   o f   S y m b o l s  S i z e   o f   O p t i o n a l   H e a d e r  C h a r a c t e r i s t i c s  M a g i c  L i n k e r   V e r s i o n  S i z e   o f   C o d e  S i z e   o f   I n i t i a l i z e d   D a t a    U n k n o w n   P E   t a r g e t  N o t   a   r e s o u r c e   d i r e c t o r y , F e a t u r e   i s   n o t   a v a i l a b l e   f o r   a t t a c h e d   i m a g e s  S e c t i o n   " % s "   n o t   f o u n d  E x p o r t s  I m p o r t s 	 R e s o u r c e s 
 E x c e p t i o n s  S e c u r i t y  B a s e   R e l o c a t i o n s  D e b u g  D e s c r i p t i o n  M a c h i n e   V a l u e  T L S  L o a d   c o n f i g u r a t i o n  B o u n d   I m p o r t ( F a i l e d   t o   g e t   A N S I   r e p l a c e m e n t   c h a r a c t e r % T h i s   W i n d o w s   v e r s i o n   i s   n o t   s u p p o r t e d & T h e   w i n d o w   w i t h   h a n d l e   % d   i s   n o t   v a l i d # T h e   p r o c e s s   w i t h   I D   % d   i s   n o t   v a l i d & T h e   m o d u l e   w i t h   h a n d l e   % d   i s   n o t   v a l i d $ F i l e   c o n t a i n s   n o   v e r s i o n   i n f o r m a t i o n  T h e   f i l e   % s   d o e s   n o t   e x i s t  I l l e g a l   l a n g u a g e   i n d e x  N o   v a l u e   w a s   s u p p l i e d  T h e   v a l u e   % s   w a s   n o t   f o u n d .  F a i l e d   t o   c r e a t e   F i l e M a p p i n g   F a i l e d   t o   c r e a t e   F i l e M a p p i n g V i e w  F a i l e d   t o   o b t a i n   s i z e   o f   f i l e  S t r e a m   i s   r e a d - o n l y  C a n n o t   o p e n   f i l e   " % s "  T h i s   i s   n o t   a   P E   f o r m a t d T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   a n   u n k n o w n   c r i t i c a l   p a r t   w h i c h   c o u l d   n o t   b e   d e c o d e d . p T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   e n c o d e d   w i t h   a n   u n k n o w n   c o m p r e s s i o n   s c h e m e   w h i c h   c o u l d   n o t   b e   d e c o d e d . c T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   u s e s   a n   u n k n o w n   i n t e r l a c e   s c h e m e   w h i c h   c o u l d   n o t   b e   d e c o d e d . ] T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   u s e s   a n   u n k n o w n   c o l o r   t y p e   w h i c h   c o u l d   n o t   b e   d e c o d e d . - T h e   c h u n k s   m u s t   b e   c o m p a t i b l e   t o   b e   a s s i g n e d . j T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   i n v a l i d   b e c a u s e   t h e   d e c o d e r   f o u n d   a n   u n e x p e c t e d   e n d   o f   t h e   f i l e . 8 T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   n o   d a t a . ] T h e   p r o g r a m   t r i e d   t o   a d d   a   e x i s t e n t   c r i t i c a l   c h u n k   t o   t h e   c u r r e n t   i m a g e   w h i c h   i s   n o t   a l l o w e d . I I t ' s   n o t   a l l o w e d   t o   a d d   a   n e w   c h u n k   b e c a u s e   t h e   c u r r e n t   i m a g e   i s   i n v a l i d . 7 T h e   p n g   i m a g e   c o u l d   n o t   b e   l o a d e d   f r o m   t h e   r e s o u r c e   I D . o S o m e   o p e r a t i o n   c o u l d   n o t   b e   p e r f o r m e d   b e c a u s e   t h e   s y s t e m   i s   o u t   o f   r e s o u r c e s .   C l o s e   s o m e   w i n d o w s   a n d   t r y   a g a i n . � S e t t i n g   b i t   t r a n s p a r e n c y   c o l o r   i s   n o t   a l l o w e d   f o r   p n g   i m a g e s   c o n t a i n i n g   a l p h a   v a l u e   f o r   e a c h   p i x e l   ( C O L O R _ R G B A L P H A   a n d   C O L O R _ G R A Y S C A L E A L P H A ) O T h i s   o p e r a t i o n   i s   n o t   v a l i d   b e c a u s e   t h e   c u r r e n t   i m a g e   c o n t a i n s   n o   v a l i d   h e a d e r . 4 T h e   n e w   s i z e   p r o v i d e d   f o r   i m a g e   r e s i z i n g   i s   i n v a l i d . o T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   c o u l d   n o t   b e   c r e a t e d   b e c a u s e   i n v a l i d   i m a g e   t y p e   p a r a m e t e r s   h a v e   b e i n g   p r o v i d e d . e T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o u l d   n o t   b e   l o a d e d   b e c a u s e   i t   u s e s   a n   i n v a l i d   i m a g e   b i t   d e p t h . 0 E l e m e n t   " % s "   d o e s   n o t   c o n t a i n   a   s i n g l e   t e x t   n o d e 4 D O M   I m p l e m e n t a t i o n   d o e s   n o t   s u p p o r t   I D O M P a r s e O p t i o n s # I t e m T a g   p r o p e r t y   i s   n o t   i n i t i a l i z e d  N o d e   i s   r e a d o n l y C R e f r e s h   i s   o n l y   s u p p o r t e d   i f   t h e   F i l e N a m e   o r   X M L   p r o p e r t i e s   a r e   s e t  F i l e N a m e   c a n n o t   b e   b l a n k  L i n e j T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   v a l i d   b e c a u s e   i t   c o n t a i n s   i n v a l i d   p i e c e s   o f   d a t a   ( c r c   e r r o r ) y T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o u l d   n o t   b e   l o a d e d   b e c a u s e   o n e   o f   i t s   m a i n   p i e c e   o f   d a t a   ( i h d r )   m i g h t   b e   c o r r u p t e d U T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   i n v a l i d   b e c a u s e   i t   h a s   m i s s i n g   i m a g e   p a r t s . [ C o u l d   n o t   d e c o m p r e s s   t h e   i m a g e   b e c a u s e   i t   c o n t a i n s   i n v a l i d   c o m p r e s s e d   d a t a .  
   D e s c r i p t i o n :   B T h e   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   c o n t a i n s   a n   i n v a l i d   p a l e t t e . � T h e   f i l e   b e i n g   r e a d   i s   n o t   a   v a l i d   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   b e c a u s e   i t   c o n t a i n s   a n   i n v a l i d   h e a d e r .   T h i s   f i l e   m a y   b e   c o r r u p t e d ,   t r y   o b t a i n i n g   i t   a g a i n n T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   s u p p o r t e d   o r   i t   m i g h t   b e   i n v a l i d .  
 ( I H D R   c h u n k   i s   n o t   t h e   f i r s t ) � T h i s   " P o r t a b l e   N e t w o r k   G r a p h i c s "   i m a g e   i s   n o t   s u p p o r t e d   b e c a u s e   e i t h e r   i t s   w i d t h   o r   h e i g h t   e x c e e d s   t h e   m a x i m u m   s i z e   o f   6 5 5 3 5   p i x e l s .  T h e r e   i s   n o   s u c h   p a l e t t e   e n t r y . C C a n n o t   c h a n g e   P o s i t i o n   o f   a   T T B D o c k   i f   i t   a l r e a d y   c o n t a i n s   c o n t r o l s G C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   N a m e   p r o p e r t y   i s   n o t   s e t O C a n n o t   s a v e   d o c k a b l e   w i n d o w ' s   p o s i t i o n   b e c a u s e   D o c k e d T o ' s   N a m e   p r o p e r t y   n o t   s e t ) " % s "   D O M I m p l e m e n t a t i o n   a l r e a d y   r e g i s t e r e d  N o   m a t c h i n g   D O M   V e n d o r :   " % s " < S e l e c t e d   D O M   V e n d o r   d o e s   n o t   s u p p o r t   t h i s   p r o p e r t y   o r   m e t h o d ; P r o p e r t y   o r   M e t h o d   " % s "   i s   n o t   s u p p o r t e d   b y   D O M   V e n d o r   " % s "  N o   s e l e c t e d   D O M   V e n d o r  N o d e   c a n n o t   b e   n u l l   M i c r o s o f t   M S X M L   i s   n o t   i n s t a l l e d  N o   a c t i v e   d o c u m e n t  N o d e   " % s "   n o t   f o u n d  I D O M N o d e   r e q u i r e d . A t t r i b u t e s   a r e   n o t   s u p p o r t e d   o n   t h i s   n o d e   t y p e  I n v a l i d   n o d e   t y p e + M i s m a t c h e d   p a r a m a t e r s   t o   R e g i s t e r C h i l d N o d e s  E x t  % s   � r   e n   o g i l t i g   e n h e t s b o k s t a v .  R � t t i g h e t e r  � g a r e  G r u p p  M � l   l � n k  F i l t y p  & K o p i e r a   h i t  & F l y t t a   h i t  & S k a p a   g e n v � g   h i t  & A v b r y t  T o o l b a r   i t e m   i n d e x   o u t   o f   r a n g e  T o o l b a r   i t e m   a l r e a d y   i n s e r t e d ? A n   i t e m   v i e w e r   a s s o c i a t e d   t h e   s p e c i f i e d   i t e m   c o u l d   n o t   b e   f o u n d  M o r e   B u t t o n s | J A   T T B D o c k   c o n t r o l   c a n n o t   b e   p l a c e d   i n s i d e   a   t o o l   w i n d o w   o r   a n o t h e r   T T B D o c k ) K a n   i n t e   b y t a   n a m n   p �   f i l   e l l e r   k a t a l o g :    F i l e n   f i n n s   r e d a n :   % F i l n a m n e t   i n n e h � l l e r   o g i l t i g a   t e c k e n :  F i l   % s  % u   F i l e r  % u   K a t a l o g e r  H u v u d k a t a l o g  D r a g D r o p   E r r o r :   % d  E n h e t   ' % s : '   � r   i n t e   k l a r .  K a t a l o g e n   ' % s '   f i n n s   i n t e .  /   < r o o t >  N a m n  S t o r l e k  F i l t y p  � n d r a d  A t t r   $ F a i l e d   t o   s e t   c a l e n d a r   m i n / m a x   r a n g e % F a i l e d   t o   s e t   c a l e n d a r   s e l e c t e d   r a n g e " ' % s '   i s   n o t   a   v a l i d   p r o p e r t y   v a l u e  O L E   c o n t r o l   a c t i v a t i o n   f a i l e d * C o u l d   n o t   o b t a i n   O L E   c o n t r o l   w i n d o w   h a n d l e % L i c e n s e   i n f o r m a t i o n   f o r   % s   i s   i n v a l i d P L i c e n s e   i n f o r m a t i o n   f o r   % s   n o t   f o u n d .   Y o u   c a n n o t   u s e   t h i s   c o n t r o l   i n   d e s i g n   m o d e N U n a b l e   t o   r e t r i e v e   a   p o i n t e r   t o   a   r u n n i n g   o b j e c t   r e g i s t e r e d   w i t h   O L E   f o r   % s / % s  B l � d d r a  A l l a   f i l e r   ( * . * ) | * . *  O g i l t i g t   f i l n a m n   -   % s # K a n   i n t e   h i t t a   n � g o n   g i l t i g   s � k v � g .  B  K B  M B  G B    I n v a l i d   i t e m   l e v e l   a s s i g n m e n t   I n v a l i d   l e v e l   ( % d )   f o r   i t e m   " % s "  I n v a l i d   i n d e x  U n a b l e   t o   i n s e r t   a n   i t e m  I n v a l i d   o w n e r  R i c h E d i t   l i n e   i n s e r t i o n   e r r o r  F a i l e d   t o   L o a d   S t r e a m  F a i l e d   t o   S a v e   S t r e a m   % s   i s   a l r e a d y   a s s o c i a t e d   w i t h   % s E % d   i s   a n   i n v a l i d   P a g e I n d e x   v a l u e .     P a g e I n d e x   m u s t   b e   b e t w e e n   0   a n d   % d = T h i s   c o n t r o l   r e q u i r e s   v e r s i o n   4 . 7 0   o r   g r e a t e r   o f   C O M C T L 3 2 . D L L  D a t e   e x c e e d s   m a x i m u m   o f   % s  D a t e   i s   l e s s   t h a n   m i n i m u m   o f   % s 4 Y o u   m u s t   b e   i n   S h o w C h e c k b o x   m o d e   t o   s e t   t o   t h i s   d a t e # F a i l e d   t o   s e t   c a l e n d a r   d a t e   o r   t i m e % F a i l e d   t o   s e t   m a x i m u m   s e l e c t i o n   r a n g e    I n v a l i d   s t y l e   f o r m a t ) C l a s s   ' % s '   i s   a l r e a d y   r e g i s t e r e d   f o r   ' % s ' % C l a s s   ' % s '   i s   n o t   r e g i s t e r e d   f o r   ' % s '  % s   p a r a m e t e r   c a n n o t   b e   n i l # F e a t u r e   n o t   s u p p o r t e d   b y   t h i s   s t y l e  S t y l e   ' % s '   i s   n o t   r e g i s t e r e d " C a n n o t   u n r e g i s t e r   t h e   s y s t e m   s t y l e  S t y l e   n o t   r e g i s t e r e d D C a n n o t   c a l l   B e g i n I n v o k e   o n   a   c o n t r o l   w i t h   n o   p a r e n t   o r   w i n d o w   h a n d l e  F a i l e d   t o   c l e a r   t a b   c o n t r o l   F a i l e d   t o   d e l e t e   t a b   a t   i n d e x   % d " F a i l e d   t o   r e t r i e v e   t a b   a t   i n d e x   % d   F a i l e d   t o   g e t   o b j e c t   a t   i n d e x   % d " F a i l e d   t o   s e t   t a b   " % s "   a t   i n d e x   % d   F a i l e d   t o   s e t   o b j e c t   a t   i n d e x   % d < M u l t i L i n e   m u s t   b e   T r u e   w h e n   T a b P o s i t i o n   i s   t p L e f t   o r   t p R i g h t % C a n n o t   r e m o v e   s h e l l   n o t i f i c a t i o n   i c o n " P a g e C o n t r o l   m u s t   f i r s t   b e   a s s i g n e d " % s   r e q u i r e s   W i n d o w s   V i s t a   o r   l a t e r  B u t t o n % d  R a d i o B u t t o n % d  C a p t i o n   c a n n o t   b e   e m p t y : C a t e g o r y P a n e l   m u s t   h a v e   a   C a t e g o r y P a n e l G r o u p   a s   i t s   p a r e n t = O n l y   C a t e g o r y P a n e l s   c a n   b e   i n s e r t e d   i n t o   a   C a t e g o r y P a n e l G r o u p  N o   h e l p   k e y w o r d   s p e c i f i e d .  U n a b l e   t o   l o a d   s t y l e   ' % s '  U n a b l e   t o   l o a d   s t y l e s :   % s  S t y l e   ' % s '   a l r e a d y   r e g i s t e r e d # S t y l e   c l a s s   ' % s '   a l r e a d y   r e g i s t e r e d  S t y l e   ' % s '   n o t   f o u n d  S t y l e   c l a s s   ' % s '   n o t   f o u n d  I n v a l i d   s t y l e   h a n d l e  P r o m p t   a r r a y   m u s t   n o t   b e   e m p t y 	 & U s e r n a m e 	 & P a s s w o r d  & D o m a i n  L o g i n 	 S e p a r a t o r  E r r o r   s e t t i n g   % s . C o u n t 8 L i s t b o x   ( % s )   s t y l e   m u s t   b e   v i r t u a l   i n   o r d e r   t o   s e t   C o u n t # N o   O n G e t I t e m   e v e n t   h a n d l e r   a s s i g n e d  " % s "   i s   a n   i n v a l i d   p a t h  A N S I  A S C I I  U n i c o d e  B i g   E n d i a n   U n i c o d e  U T F - 8  U T F - 7     C l i p b o a r d   d o e s   n o t   s u p p o r t   I c o n s  C a n n o t   o p e n   c l i p b o a r d :   % s  T e x t   e x c e e d s   m e m o   c a p a c i t y + O p e r a t i o n   n o t   s u p p o r t e d   o n   s e l e c t e d   p r i n t e r . T h e r e   i s   n o   d e f a u l t   p r i n t e r   c u r r e n t l y   s e l e c t e d / M e n u   ' % s '   i s   a l r e a d y   b e i n g   u s e d   b y   a n o t h e r   f o r m  P i c t u r e :    ( % d x % d )  P r e v i e w  D o c k e d   c o n t r o l   m u s t   h a v e   a   n a m e % E r r o r   r e m o v i n g   c o n t r o l   f r o m   d o c k   t r e e    -   D o c k   z o n e   n o t   f o u n d    -   D o c k   z o n e   h a s   n o   c o n t r o l L E r r o r   l o a d i n g   d o c k   z o n e   f r o m   t h e   s t r e a m .   E x p e c t i n g   v e r s i o n   % d ,   b u t   f o u n d   % d . , M u l t i s e l e c t   m o d e   m u s t   b e   o n   f o r   t h i s   f e a t u r e 7 L e n g t h   o f   v a l u e   a r r a y   m u s t   b e   > =   l e n g t h   o f   p r o m p t   a r r a y  E n d  H o m e  L e f t  U p  R i g h t  D o w n  I n s  D e l  S h i f t +  C t r l +  A l t +  ( N o n e )  V a l u e   m u s t   b e   b e t w e e n   % d   a n d   % d  A l l  U n a b l e   t o   i n s e r t   a   l i n e  I n v a l i d   c l i p b o a r d   f o r m a t  A v b r y t  & H j � l p  & A v b r y t  & F � r s � k   i g e n 	 & I g n o r e r a  & A l l a  N & e j   t i l l   a l l a  J & a   t i l l   a l l a  & S t � n g  B k S p  T a b  E s c  E n t e r  S p a c e  P g U p  P g D n  T I F F   I m a g e s  G r i d   t o o   l a r g e   f o r   o p e r a t i o n   T o o   m a n y   r o w s   o r   c o l u m n s   d e l e t e d  G r i d   i n d e x   o u t   o f   r a n g e 1 F i x e d   c o l u m n   c o u n t   m u s t   b e   l e s s   t h a n   c o l u m n   c o u n t + F i x e d   r o w   c o u n t   m u s t   b e   l e s s   t h a n   r o w   c o u n t & C a n n o t   i n s e r t   o r   d e l e t e   r o w s   f r o m   g r i d  O g i l t i g t   i n p u t v � r d e 9 O g i l t i g t   i n p u t v � r d e .   A n v � n d   E S C   f � r   a t t   a v b r y t a   � n d r i n g a r  V a r n i n g  F e l  I n f o r m a t i o n  B e k r � f t a  & J a  & N e j  O K ) C o n t r o l   ' % s '   i s   u s e d   o n   a   n o t   m a i n   t h r e a d  O K  A v b r y t  & Y e s  & N o  & H e l p  & C l o s e  & I g n o r e  & R e t r y  A b o r t  & A l l  C a n n o t   d r a g   a   f o r m 	 M e t a f i l e s  E n h a n c e d   M e t a f i l e s  I c o n s  B i t m a p s  % s   p r o p e r t y   o u t   o f   r a n g e 3 C h e c k   s t a t e   c a n   o n l y   b e   s e t   w h e n   C h e c k B o x e s   i s   T r u e 4 C h e c k   s t a t e   i n c o m p a t i b l e   w i t h   t r e e v i e w ' s   C h e c k S t y l e s  M e n u   i n d e x   o u t   o f   r a n g e  M e n u   i n s e r t e d   t w i c e  S u b - m e n u   i s   n o t   i n   m e n u  N o t   e n o u g h   t i m e r s   a v a i l a b l e ! P r i n t e r   i s   n o t   c u r r e n t l y   p r i n t i n g  P r i n t i n g   i n   p r o g r e s s  P r i n t e r   i n d e x   o u t   o f   r a n g e  P r i n t e r   s e l e c t e d   i s   n o t   v a l i d  % s   o n   % s @ G r o u p I n d e x   c a n n o t   b e   l e s s   t h a n   a   p r e v i o u s   m e n u   i t e m ' s   G r o u p I n d e x 5 C a n n o t   c r e a t e   f o r m .   N o   M D I   f o r m s   a r e   c u r r e n t l y   a c t i v e 0 C a n   o n l y   m o d i f y   a n   i m a g e   i f   i t   c o n t a i n s   a   b i t m a p * A   c o n t r o l   c a n n o t   h a v e   i t s e l f   a s   i t s   p a r e n t  I n v a l i d   I m a g e L i s t  U n a b l e   t o   R e p l a c e   I m a g e  U n a b l e   t o   I n s e r t   I m a g e  I n v a l i d   I m a g e L i s t   I n d e x ) F a i l e d   t o   r e a d   I m a g e L i s t   d a t a   f r o m   s t r e a m ( F a i l e d   t o   w r i t e   I m a g e L i s t   d a t a   t o   s t r e a m $ E r r o r   c r e a t i n g   w i n d o w   d e v i c e   c o n t e x t  E r r o r   c r e a t i n g   w i n d o w   c l a s s + C a n n o t   f o c u s   a   d i s a b l e d   o r   i n v i s i b l e   w i n d o w ! C o n t r o l   ' % s '   h a s   n o   p a r e n t   w i n d o w  .   P a t h :  
 % s $ P a r e n t   g i v e n   i s   n o t   a   p a r e n t   o f   ' % s '  C a n n o t   h i d e   a n   M D I   C h i l d   F o r m ) C a n n o t   c h a n g e   V i s i b l e   i n   O n S h o w   o r   O n H i d e " C a n n o t   m a k e   a   v i s i b l e   w i n d o w   m o d a l  S c r o l l b a r   p r o p e r t y   o u t   o f   r a n g e    I c o n   i m a g e   i s   n o t   v a l i d  M e t a f i l e   i s   n o t   v a l i d  I n v a l i d   p i x e l   f o r m a t  I n v a l i d   i m a g e  S c a n   l i n e   i n d e x   o u t   o f   r a n g e ! C a n n o t   c h a n g e   t h e   s i z e   o f   a n   i c o n % C a n n o t   c h a n g e   t h e   s i z e   o f   a   W I C   I m a g e   I n v a l i d   o p e r a t i o n   o n   T O l e G r a p h i c $ U n k n o w n   p i c t u r e   f i l e   e x t e n s i o n   ( . % s )  U n s u p p o r t e d   c l i p b o a r d   f o r m a t  U n s u p p o r t e d   s t r e a m   f o r m a t  O u t   o f   s y s t e m   r e s o u r c e s  C a n v a s   d o e s   n o t   a l l o w   d r a w i n g # T e x t   f o r m a t   f l a g   ' % s '   n o t   s u p p o r t e d 8 I n v a l i d   i m a g e   f r a m e   i n d e x   % d :   t h e r e   a r e   % d   f r a m e s   ( 0 - % d )  I n v a l i d   i m a g e   s i z e    E r r o r   r e a d i n g   d a t a :   ( % d )   % s . E r r o r   s e t t i n g   t i m e o u t   f o r   t h e   r e q u e s t :   ( % d )   % s ' E r r o r   o p e n i n g   c e r t i f i c a t e   f i l e :   ( % d )   % s ) C e r t i f i c a t e   i s   n o t   f o u n d   i n   f i l e :   ( % d )   % s . P a i r   o f   e x t e n s i o n   a n d   m i m e   t y p e   a l r e a d y   e x i s t s  M i m e   t y p e   c a n n o t   b e   e m p t y  V a l u e   n a m e   c a n n o t   b e   e m p t y  Q u a l i t y   w e i g h t   i s   o u t   o f   r a n g e  O L E   e r r o r   % . 8 x . M e t h o d   ' % s '   n o t   s u p p o r t e d   b y   a u t o m a t i o n   o b j e c t / V a r i a n t   d o e s   n o t   r e f e r e n c e   a n   a u t o m a t i o n   o b j e c t 7 D i s p a t c h   m e t h o d s   d o   n o t   s u p p o r t   m o r e   t h a n   6 4   p a r a m e t e r s  D C O M   n o t   i n s t a l l e d 0 T a b   p o s i t i o n   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   s t y l e 0 T a b   s t y l e   i n c o m p a t i b l e   w i t h   c u r r e n t   t a b   p o s i t i o n  B i t m a p   i m a g e   i s   n o t   v a l i d   , M a x i m u m   n u m b e r   o f   r e d i r e c t i o n s   ( % d )   e x c e e d e d   E r r o r   g e t t i n g   S e r v e r   C e r t i f i c a t e ) S e r v e r   C e r t i f i c a t e   I n v a l i d   o r   n o t   p r e s e n t  S e r v e r   C e r t i f i c a t e   n o t   a c c e p t e d  E m p t y   c e r t i f i c a t e   l i s t # U n s p e c i f i e d   c e r t i f i c a t e   f r o m   c l i e n t  C l i e n t   r e j e c t e d   t h e   c e r t i f i c a t e 2 E x e c u t i o n   o f   r e q u e s t   t e r m i n a t e d   w i t h   u n k n o w n   e r r o r  E r r o r   q u e r y i n g   h e a d e r s :   ( % d )   % s  E r r o r   o b t a i n i n g   s e s s i o n   h a n d l e  E r r o r   s e n d i n g   d a t a :   ( % d )   % s  E r r o r   r e c e i v i n g   d a t a :   ( % d )   % s  E r r o r   c o n n e c t i n g   t o   s e r v e r :   % s  E r r o r   o p e n i n g   r e q u e s t :   ( % d )   % s  E r r o r   a d d i n g   h e a d e r :   ( % d )   % s  E r r o r   r e m o v i n g   h e a d e r :   ( % d )   % s    P a t h   e n d e d   w i t h   a n   o p e n   b r a c k e t  P a t h   e n d e d   w i t h   a n   o p e n   s t r i n g  I n v a l i d   i n d e x   f o r   a r r a y :   % s . U n e x p e c t e d   c h a r a c t e r   w h i l e   p a r s i n g   i n d e x e r :   % s 0 E m p t y   n a m e   n o t   a l l o w e d   i n   d o t   n o t a t i o n ,   u s e   [ ' ' ] % S c h e m e   " % s "   a l r e a d y   r e g i s t e r e d   f o r   % s  S c h e m e   " % s "   i s   n o t   r e g i s t e r e d $ C r e d e n t i a l   w i t h o u t   u s e r   a n d   p a s s w o r d + P l a t f o r m - d e p e n d a n t   f u n c t i o n   n o t   i m p l e m e n t e d ) S c h e m e - d e p e n d a n t   f u n c t i o n   n o t   i m p l e m e n t e d  M e t h o d   a l r e a d y   a s s i g n e d  U R L   a l r e a d y   a s s i g n e d * P a r a m e t e r   i n d e x   ( % d )   o u t   o f   r a n g e   ( % d . . % d )  I n v a l i d   U R L :   " % s "  P a r a m e t e r   " % s "   n o t   f o u n d  I n v a l i d   r e l a t i v e   U R L   p a t h :   " % s "    N o   t o k e n   t o   c l o s e . . T h e   r e a d e r ' s   M a x D e p t h   o f   % s   h a s   b e e n   e x c e e d e d . < T o k e n   % s   i n   s t a t e   % s   w o u l d   r e s u l t   i n   a n   i n v a l i d   J S O N   o b j e c t . " U n e x p e c t e d   e n d   w h e n   r e a d i n g   b y t e s . , U n e x p e c t e d   e n d   w h e n   r e a d i n g   d a t e   c o n s t r u c t o r ( E r r o r   r e a d i n g   d a t e .   U n e x p e c t e d   t o k e n :   % s O U n e x p e c t e d   t o k e n   w h e n   r e a d i n g   d a t e   c o n s t r u c t o r .   E x p e c t e d   E n d C o n s t r u c t o r ,   g o t   % s H U n e x p e c t e d   t o k e n   w h e n   r e a d i n g   d a t e   c o n s t r u c t o r .   E x p e c t e d   I n t e g e r ,   g o t   % s * E r r o r   r e a d i n g   d o u b l e .   U n e x p e c t e d   t o k e n :   % s + E r r o r   r e a d i n g   i n t e g e r .   U n e x p e c t e d   t o k e n :   % s ' U n e x p e c t e d   t o k e n   w h e n   r e a d i n g   b y t e s :   % s * E r r o r   r e a d i n g   s t r i n g .   U n e x p e c t e d   t o k e n :   % s $ U n e x p e c t e d   t y p e   w h e n   w r i t i n g   e n d :   % s  U n k n o w n   J s o n T y p e :   % s  U n s u p p o r t e d   t y p e :   % s # U n e x p e c t e d   c h a r   f o r   r o o t   e l e m e n t :   . 2 U T F 8 :   T y p e   c a n n o t   b e   d e t e r m i n e d   o u t   o f   h e a d e r   b y t e # T h e   i n p u t   v a l u e   i s   n o t   a   v a l i d   J S O N - .   P a t h   ' % s ' ,   l i n e   % d ,   p o s i t i o n   % d   ( o f f s e t   % d ) = T h e   n e s t i n g   l e v e l   o f   J S O N   a r r a y s   /   o b j e c t s   i s   g r e a t e r   t h a n   % d  V a l u e   ' % s '   n o t   f o u n d  V a l u e   % s   c a n n o t   b e   a d d e d   t o   % s ( C o u l d   n o t   c o n v e r t   s t r i n g   t o   D a t e T i m e :   % s & C o u l d   n o t   c o n v e r t   s t r i n g   t o   d o u b l e :   % s ' C o u l d   n o t   c o n v e r t   s t r i n g   t o   i n t e g e r :   % s  ,   l i n e   % d ,   p o s i t i o n   % d 	 P a t h   ' % s '  N o t   a   v a l i d   c l o s e   J s o n T o k e n :   % s  A n   O b j e c t I d   m u s t   b e   1 2   b y t e s  I n v a l i d   s t a t e :   % s 2 J s o n T o k e n   % s   i s   n o t   v a l i d   f o r   c l o s i n g   J s o n T y p e   % s .  N o   c l o s e   t o k e n   f o r   t y p e   % s    A t   l e a s t   o n e   t a s k   i n   a r r a y   n i l . C a n n o t   s t a r t   a   t a s k   t h a t   h a s   a l r e a d y   c o m p l e t e d   O n e   o r   m o r e   t a s k s   w e r e   c a n c e l l e d  O n e   o r   m o r e   e r r o r s   o c c u r r e d  M u s t   w a i t   o n   a t   l e a s t   o n e   e v e n t E C a n n o t   c a l l   B e g i n I n v o k e   o n   a   T C o m p o n e n t   i n   t h e   p r o c e s s   o f   d e s t r u c t i o n 3 A   r e g u l a r   e x p r e s s i o n   s p e c i f i e d   i n   R e g E x   i s   r e q u i r e d , E r r o r   i n   r e g u l a r   e x p r e s s i o n   a t   o f f s e t   % d :   % s  E r r o r   s t u d y i n g   t h e   r e g e x :   % s  S u c c e s s f u l   m a t c h   r e q u i r e d  S t r i n g s   p a r a m e t e r   c a n n o t   b e   n i l  I n v a l i d   i n d e x   t y p e  I n d e x   o u t   o f   b o u n d s   ( % d )  I n v a l i d   g r o u p   n a m e   ( % s ) < U T F 8 :   A   s t a r t   b y t e   n o t   f o l l o w e d   b y   e n o u g h   c o n t i n u a t i o n   b y t e s 5 U T F 8 :   A n   u n e x p e c t e d   c o n t i n u a t i o n   b y t e   i n   % d - b y t e   U T F 8 
 W i n d o w s   1 0 
 W i n d o w s   1 1 " C a n n o t   c r e a t e   i n s t a n c e   o f   c l a s s   % s  O b s e r v e r   i s   n o t   s u p p o r t e d L C a n n o t   h a v e   m u l t i p l e   s i n g l e   c a s t   o b s e r v e r s   a d d e d   t o   t h e   o b s e r v e r s   c o l l e c t i o n 4 T h e   o b j e c t   d o e s   n o t   i m p l e m e n t   t h e   o b s e r v e r   i n t e r f a c e G N o   s i n g l e   c a s t   o b s e r v e r   w i t h   I D   % d   w a s   a d d e d   t o   t h e   o b s e r v e r   c o l l e c t i o n F N o   m u l t i   c a s t   o b s e r v e r   w i t h   I D   % d   w a s   a d d e d   t o   t h e   o b s e r v e r   c o l l e c t i o n  O b s e r v e r   i s   n o t   a v a i l a b l e  I n v a l i d   d a t e   s t r i n g :   % s  I n v a l i d   t i m e   s t r i n g :   % s  I n v a l i d   t i m e   O f f s e t   s t r i n g :   % s = E r r o r   d e c o d i n g   U R L   s t y l e   ( % % X X )   e n c o d e d   s t r i n g   a t   p o s i t i o n   % d 1 I n v a l i d   U R L   e n c o d e d   c h a r a c t e r   ( % s )   a t   p o s i t i o n   % d ( C a n n o t   c o n s t r u c t   a n   I T a s k   i n   t h i s   m a n n e r " L i s t   o f   t a s k s   t o   J o i n   m e t h o d   e m p t y    W i n d o w s  W i n d o w s   V i s t a  W i n d o w s   S e r v e r   2 0 0 8 	 W i n d o w s   7  W i n d o w s   S e r v e r   2 0 0 8   R 2  W i n d o w s   2 0 0 0 
 W i n d o w s   X P  W i n d o w s   S e r v e r   2 0 0 3  W i n d o w s   S e r v e r   2 0 0 3   R 2  W i n d o w s   S e r v e r   2 0 1 2  W i n d o w s   S e r v e r   2 0 1 2   R 2  W i n d o w s   S e r v e r   2 0 1 6  W i n d o w s   S e r v e r   2 0 1 9  W i n d o w s   S e r v e r   2 0 2 2 	 W i n d o w s   8  W i n d o w s   8 . 1    A r g u m e n t   m u s t   n o t   b e   n i l # U n b a l a n c e d   s t a c k   o r   q u e u e   o p e r a t i o n  I t e m   n o t   f o u n d  D u p l i c a t e s   n o t   a l l o w e d  T h r e a d   t r a c k i n g   i s n ' t   e n a b l e d / S p i n L o c k   h a s   b e e n   r e - e n t e r e d   o n   t h e   s a m e   t h r e a d ( S p i n L o c k   n o t   o w n e d   b y   t h e   c u r r e n t   t h r e a d 5 I n s u f f i c i e n t   R T T I   a v a i l a b l e   t o   s u p p o r t   t h i s   o p e r a t i o n  P a r a m e t e r   c o u n t   m i s m a t c h < T y p e   ' % s '   i s   n o t   d e c l a r e d   i n   t h e   i n t e r f a c e   s e c t i o n   o f   a   u n i t 7 V A R   a n d   O U T   a r g u m e n t s   m u s t   m a t c h   p a r a m e t e r   t y p e   e x a c t l y , S p e c i f i e d   L o g i n   C r e d e n t i a l   S e r v i c e   n o t   f o u n d " % s   ( V e r s i o n   % d . % d ,   B u i l d   % d ,   % 5 : s ) : % s   S e r v i c e   P a c k   % 4 : d   ( V e r s i o n   % 1 : d . % 2 : d ,   B u i l d   % 3 : d ,   % 5 : s )  3 2 - b i t   E d i t i o n  6 4 - b i t   E d i t i o n   + C o u n t   a l r e a d y   m a x :   A m o u n t :   % d ,   C u r C o u n t :   % d " C o u n t d o w n   a l r e a d y   r e a c h e d   z e r o   ( 0 )  T i m e s p a n   t o o   l o n g b T h e   d u r a t i o n   c a n n o t   b e   r e t u r n e d   b e c a u s e   t h e   a b s o l u t e   v a l u e   e x c e e d s   t h e   v a l u e   o f   T T i m e S p a n . M a x V a l u e  V a l u e   c a n n o t   b e   N a N 3 N e g a t i n g   t h e   m i n i m u m   v a l u e   o f   a   T i m e s p a n   i s   i n v a l i d  I n v a l i d   T i m e s p a n   f o r m a t  T i m e s p a n   e l e m e n t   t o o   l o n g # N o   c o n t e x t - s e n s i t i v e   h e l p   i n s t a l l e d  N o   h e l p   f o u n d   f o r   c o n t e x t   % d  U n a b l e   t o   o p e n   I n d e x  U n a b l e   t o   o p e n   S e a r c h " U n a b l e   t o   f i n d   a   T a b l e   o f   C o n t e n t s $ N o   t o p i c - b a s e d   h e l p   s y s t e m   i n s t a l l e d  N o   h e l p   f o u n d   f o r   % s  A r g u m e n t   o u t   o f   r a n g e   , ( % d ,   % d ,   % d )   i s   n o t   a   v a l i d   D a t e W e e k   t r i p l e t  ? W T h e   g i v e n   " % s "   l o c a l   t i m e   i s   i n v a l i d   ( s i t u a t e d   w i t h i n   t h e   m i s s i n g   p e r i o d   p r i o r   t o   D S T ) . $ N o   h e l p   v i e w e r   t h a t   s u p p o r t s   f i l t e r s  I n v a l i d   a r g u m e n t / I n d e x   o u t   o f   r a n g e   ( % d ) .     M u s t   b e   > =   0   a n d   <   % d 2 L e n g t h   o f   S t r i n g s   a n d   O b j e c t s   a r r a y s   m u s t   b e   e q u a l 2 S o u r c e   a n d   D e s t i n a t i o n   a r r a y s   m u s t   n o t   b e   t h e   s a m e * C l a s s   % s   i s   n o t   i n t e n d e d   t o   b e   c o n s t r u c t e d  I n v a l i d   T i m e o u t   v a l u e :   % s 0 S p i n C o u n t   o u t   o f   r a n g e .   M u s t   b e   b e t w e e n   0   a n d   % d  I n v a l i d   R e s e t   C o u n t :   % d  I n v a l i d   C o u n t :   % d  I n v a l i d   D e c r e m e n t   C o u n t :   % d  I n v a l i d   I n c r e m e n t   C o u n t :   % d D D e c r e m e n t   a m o u n t   w i l l   c a u s e   i n v a l i d   r e s u l t s :   C o u n t :   % d ,   C u r C o u n t :   % d 9 C a n n o t   c a l l   S e t R e t u r n V a l u e   o n   a n   e x t e r n a l l y   c r e a t e   t h r e a d  P a r a m e t e r   % s   c a n n o t   b e   n i l ' P a r a m e t e r   % s   c a n n o t   b e   a   n e g a t i v e   v a l u e * I n p u t   b u f f e r   e x c e e d e d   f o r   % s   =   % d ,   % s   =   % d  I n v a l i d   c h a r a c t e r s   i n   p a t h  I n v a l i d   c h a r a c t e r s   i n   f i l e   n a m e  P a t h   i s   e m p t y  F i l e   n a m e   i s   e m p t y  T h e   s p e c i f i e d   p a t h   i s   t o o   l o n g   T h e   s p e c i f i e d   p a t h   w a s   n o t   f o u n d   T h e   p a t h   f o r m a t   i s   n o t   s u p p o r t e d  T h e   d r i v e   c a n n o t   b e   f o u n d   T h e   s p e c i f i e d   f i l e   w a s   n o t   f o u n d ! T h e   s p e c i f i e d   f i l e   a l r e a d y   e x i s t s  T h e   s p e c i f i e d   f i l e   i s   t o o   l o n g . $ ( % d ,   % d )   i s   n o t   a   v a l i d   D a t e D a y   p a i r    F a i l e d   t o   c r e a t e   k e y   % s  F a i l e d   t o   g e t   d a t a   f o r   ' % s '  I n v a l i d   c o m p o n e n t   r e g i s t r a t i o n  F a i l e d   t o   s e t   d a t a   f o r   ' % s '  R e s o u r c e   % s   n o t   f o u n d  % s . S e e k   n o t   i m p l e m e n t e d $ O p e r a t i o n   n o t   a l l o w e d   o n   s o r t e d   l i s t $ % s   n o t   i n   a   c l a s s   r e g i s t r a t i o n   g r o u p  P r o p e r t y   % s   d o e s   n o t   e x i s t  S t r e a m   w r i t e   e r r o r  T h r e a d   c r e a t i o n   e r r o r :   % s  T h r e a d   E r r o r :   % s   ( % d ) - C a n n o t   t e r m i n a t e   a n   e x t e r n a l l y   c r e a t e d   t h r e a d , C a n n o t   w a i t   f o r   a n   e x t e r n a l l y   c r e a t e d   t h r e a d 2 C a n n o t   c a l l   S t a r t   o n   a   r u n n i n g   o r   s u s p e n d e d   t h r e a d ; C a n n o t   c a l l   C h e c k T e r m i n a t e d   o n   a n   e x t e r n a l l y   c r e a t e d   t h r e a d    ' % s '   i s   a n   i n v a l i d   m a s k   a t   ( % d ) $ ' ' % s ' '   i s   n o t   a   v a l i d   c o m p o n e n t   n a m e  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   p r o p e r t y   e l e m e n t :   % s  I n v a l i d   p r o p e r t y   p a t h  I n v a l i d   p r o p e r t y   t y p e :   % s  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   d a t a   t y p e   f o r   ' % s '   L i s t   c a p a c i t y   o u t   o f   b o u n d s   ( % d )  L i s t   c o u n t   o u t   o f   b o u n d s   ( % d )  L i s t   i n d e x   o u t   o f   b o u n d s   ( % d ) + O u t   o f   m e m o r y   w h i l e   e x p a n d i n g   m e m o r y   s t r e a m ) % s   h a s   n o t   b e e n   r e g i s t e r e d   a s   a   C O M   c l a s s  E r r o r   r e a d i n g   % s % s % s :   % s  S t r e a m   r e a d   e r r o r  P r o p e r t y   i s   r e a d - o n l y    I n v a l i d   S t r i n g B a s e I n d e x  O p e r a t i o n   C a n c e l l e d  A n c e s t o r   f o r   ' % s '   n o t   f o u n d  C a n n o t   a s s i g n   a   % s   t o   a   % s  B i t s   i n d e x   o u t   o f   r a n g e * C a n ' t   w r i t e   t o   a   r e a d - o n l y   r e s o u r c e   s t r e a m E C h e c k S y n c h r o n i z e   c a l l e d   f r o m   t h r e a d   $ % x ,   w h i c h   i s   N O T   t h e   m a i n   t h r e a d  C l a s s   % s   n o t   f o u n d  A   c l a s s   n a m e d   % s   a l r e a d y   e x i s t s % L i s t   d o e s   n o t   a l l o w   d u p l i c a t e s   ( $ 0 % x ) # A   c o m p o n e n t   n a m e d   % s   a l r e a d y   e x i s t s % S t r i n g   l i s t   d o e s   n o t   a l l o w   d u p l i c a t e s  C a n n o t   c r e a t e   f i l e   " % s " .   % s  C a n n o t   o p e n   f i l e   " % s " .   % s  U n a b l e   t o   w r i t e   t o   % s  I n v a l i d   s t r e a m   f o r m a t    M o n d a y  T u e s d a y 	 W e d n e s d a y  T h u r s d a y  F r i d a y  S a t u r d a y  U n a b l e   t o   c r e a t e   d i r e c t o r y  I n v a l i d   s o u r c e   a r r a y  I n v a l i d   d e s t i n a t i o n   a r r a y " C h a r a c t e r   i n d e x   o u t   o f   b o u n d s   ( % d )  S t a r t   i n d e x   o u t   o f   b o u n d s   ( % d )  I n v a l i d   c o u n t   ( % d )  I n v a l i d   d e s t i n a t i o n   i n d e x   ( % d )  I n v a l i d   c o d e   p a g e  I n v a l i d   e n c o d i n g   n a m e N N o   m a p p i n g   f o r   t h e   U n i c o d e   c h a r a c t e r   e x i s t s   i n   t h e   t a r g e t   m u l t i - b y t e   c o d e   p a g e    M a y  J u n e  J u l y  A u g u s t 	 S e p t e m b e r  O c t o b e r  N o v e m b e r  D e c e m b e r  S u n  M o n  T u e  W e d  T h u  F r i  S a t  S u n d a y  J a n  F e b  M a r  A p r  M a y  J u n  J u l  A u g  S e p  O c t  N o v  D e c  J a n u a r y  F e b r u a r y  M a r c h  A p r i l    E x t e r n a l   e x c e p t i o n   % x  A s s e r t i o n   f a i l e d  I n t e r f a c e   n o t   s u p p o r t e d  E x c e p t i o n   i n   s a f e c a l l   m e t h o d  O b j e c t   l o c k   n o t   o w n e d ( M o n i t o r   s u p p o r t   f u n c t i o n   n o t   i n i t i a l i z e d  % d   e x c e p t i o n ( s ) :  F e a t u r e   n o t   i m p l e m e n t e d   M e t h o d   c a l l e d   o n   d i s p o s e d   o b j e c t  % s   ( % s ,   l i n e   % d )  A b s t r a c t   E r r o r ? A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p   i n   m o d u l e   ' % s ' .   % s   o f   a d d r e s s   % p 2 C a n n o t   a c c e s s   p a c k a g e   i n f o r m a t i o n   f o r   p a c k a g e   ' % s '  C a n ' t   l o a d   p a c k a g e   % s .  
 % s  S y s t e m f e l .   K o d :   % d .  
 % s % s * E t t   a n r o p   t i l l   e n   O S   f u n k t i o n   m i s s l y c k a d e s  V a r i a n t   o r   s a f e   a r r a y   i s   l o c k e d  I n v a l i d   v a r i a n t   t y p e   c o n v e r s i o n  I n v a l i d   v a r i a n t   o p e r a t i o n  I n v a l i d   N U L L   v a r i a n t   o p e r a t i o n % I n v a l i d   v a r i a n t   o p e r a t i o n   ( % s % . 8 x ) 
 % s , C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   i s   o u t   o f   r a n g e / C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   a l r e a d y   u s e d   b y   % s * C u s t o m   v a r i a n t   t y p e   ( % s % . 4 x )   i s   n o t   u s a b l e 2 T o o   m a n y   c u s t o m   v a r i a n t   t y p e s   h a v e   b e e n   r e g i s t e r e d 5 C o u l d   n o t   c o n v e r t   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s ) = O v e r f l o w   w h i l e   c o n v e r t i n g   v a r i a n t   o f   t y p e   ( % s )   i n t o   t y p e   ( % s )  V a r i a n t   o v e r f l o w  I n v a l i d   a r g u m e n t  I n v a l i d   v a r i a n t   t y p e  O p e r a t i o n   n o t   s u p p o r t e d  U n e x p e c t e d   v a r i a n t   e r r o r  S t a c k   o v e r f l o w  C o n t r o l - C   h i t  P r i v i l e g e d   i n s t r u c t i o n  O p e r a t i o n   a b o r t e d ( E x c e p t i o n   % s   i n   m o d u l e   % s   a t   % p .  
 % s % s  
  A p p l i c a t i o n   E r r o r 1 F o r m a t   ' % s '   i n v a l i d   o r   i n c o m p a t i b l e   w i t h   a r g u m e n t  N o   a r g u m e n t   f o r   f o r m a t   ' % s ' " V a r i a n t   m e t h o d   c a l l s   n o t   s u p p o r t e d  R e a d  W r i t e 	 E x e c u t i o n  I n v a l i d   a c c e s s  F o r m a t   s t r i n g   t o o   l o n g $ E r r o r   c r e a t i n g   v a r i a n t   o r   s a f e   a r r a y ) V a r i a n t   o r   s a f e   a r r a y   i n d e x   o u t   o f   b o u n d s  T o o   m a n y   o p e n   f i l e s  F i l e   a c c e s s   d e n i e d  R e a d   b e y o n d   e n d   o f   f i l e 	 D i s k   f u l l  I n v a l i d   n u m e r i c   i n p u t  D i v i s i o n   b y   z e r o  R a n g e   c h e c k   e r r o r  I n t e g e r   o v e r f l o w   I n v a l i d   f l o a t i n g   p o i n t   o p e r a t i o n  F l o a t i n g   p o i n t   d i v i s i o n   b y   z e r o  F l o a t i n g   p o i n t   o v e r f l o w  F l o a t i n g   p o i n t   u n d e r f l o w  I n v a l i d   p o i n t e r   o p e r a t i o n  I n v a l i d   c l a s s   t y p e c a s t 0 A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p .   % s   o f   a d d r e s s   % p  A c c e s s   v i o l a t i o n 	 < u n k n o w n > ! ' % s '   i s   n o t   a   v a l i d   i n t e g e r   v a l u e - ' % s '   i s   n o t   a   v a l i d   i n t e g e r   v a l u e   f o r   % s   t y p e ( ' % s '   i s   n o t   a   v a l i d   f l o a t i n g   p o i n t   v a l u e  ' % s '   � r   i n g e t   g i l t i g t   d a t u m  ' % s '   � r   i n g e n   g i l t i g   t i d # ' % s '   � r   i n g e t   g i l t i g t   d a t u m   o c h   t i d   ' % d . % d '   i s   n o t   a   v a l i d   t i m e s t a m p  ' % s '   i s   n o t   a   v a l i d   G U I D   v a l u e ! ' % s '   i s   n o t   a   v a l i d   b o o l e a n   v a l u e  I n v a l i d   a r g u m e n t   t o   t i m e   e n c o d e  I n v a l i d   a r g u m e n t   t o   d a t e   e n c o d e  O u t   o f   m e m o r y  I / O   e r r o r   % d  F i l e   n o t   f o u n d  I n v a l i d   f i l e n a m e   &=O87��$B�:�TPF0TAboutDialogAboutDialogLeftuTop{HelpType	htKeywordHelpKeywordui_aboutBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	Om WinSCPClientHeightClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 
KeyPreview	PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChanged	OnKeyDownFormKeyDown
DesignSize� 
TextHeight TButtonOKButtonLeftTop�WidthPHeightAnchorsakRightakBottom Cancel	CaptionOKDefault	ModalResultTabOrder OnMouseDownOKButtonMouseDown  TButtonLicenseButtonLeft>Top�WidthPHeightAnchorsakLeftakBottom Caption
&Licens...TabOrderOnClickLicenseButtonClick  TButton
HelpButtonLeftoTop�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelPanelLeft Top Width�Height�AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder
DesignSize��  TLabelApplicationLabelLeft>TopWidth=HeightCaptionApplicationShowAccelChar  TLabelVersionLabelLeft>TopWidth� HeightCaptionVersion 2.0.0 (Build 12) XXShowAccelChar  TLabelWinSCPCopyrightLabelLeft>Top:Width� HeightCaption%   Copyright © 2000-2003 Martin PrikrylShowAccelChar  TLabelProductSpecificMessageLabelLeft>TophWidth1HeightCaption5   För att skicka in kommentarer och rapportera buggar:ShowAccelChar  TLabelLabel3Left>Top	WidtheHeightCaption   Copyright för vissa delar:ShowAccelChar  TLabelRegistrationLabelLeft>Top� Width� HeightCaptionThis product is licensed to:ShowAccelChar  	TPaintBoxIconPaintBoxLeftTopWidth0Height0OnPaintIconPaintBoxPaint  TStaticTextHomepageLabelLeft>TopLWidth� HeightCaptionhttp://XXXXXXwinscp.net/TabOrder TabStop	  TStaticTextForumUrlLabelLeft>TopzWidth� HeightCaptionhttp://XXXXwinscp.net/forum/TabOrderTabStop	  TPanelThirdPartyPanelLeft@TopWidthHeight� AnchorsakLeftakTopakRight 	BevelKindbkTile
BevelOuterbvNoneParentColor	TabOrder  TPanelRegistrationBoxLeft>Top� Width�HeightYAnchorsakLeftakTopakRight 	BevelKindbkTile
BevelOuterbvNoneParentBackgroundParentColor	TabOrder
DesignSize}U  TLabelRegistrationSubjectLabelLeftTopWidth HeightAAnchorsakLeftakTopakRight AutoSizeCaptionSomeone
Somewhere, some cityShowAccelCharWordWrap	  TLabelRegistrationLicensesLabelLeftTop+WidthvHeightCaptionNumber of Licenses: XShowAccelChar  TStaticTextRegistrationProductIdLabelLeftTopAWidth� HeightCaptionProduct ID: xxxx-xxxx-xxxxxShowAccelCharTabOrder OnClickRegistrationProductIdLabelClick        TPF0TAuthenticateFormAuthenticateFormLeft0TopqHelpType	htKeywordHelpKeywordui_authenticateBorderIconsbiSystemMenu BorderStylebsDialogCaptionAuthenticateFormClientHeight|ClientWidth�Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidthFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnResize
FormResizeOnShowFormShow
TextHeight TPanelTopPanelLeft Top Width�Height?AlignalClient
BevelOuterbvNoneTabOrder  TListBoxLogViewLeft0Top WidthpHeight?StylelbOwnerDrawVariableAlignalClient
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneDoubleBuffered	ParentDoubleBufferedParentShowHintShowHint	TabOrder 
OnDrawItemLogViewDrawItemOnMeasureItemLogViewMeasureItemOnMouseMoveLogViewMouseMove  TPanel	LeftPanelLeft Top Width0Height?AlignalLeft
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder 	TPaintBoxAnimationPaintBoxLeftTopWidth Height     TPanelPasswordPanelLeft Top?Width�Height� AlignalBottomAutoSize	
BevelOuterbvNoneTabOrderVisible TPanelPromptEditPanelLeft Top Width�Height� AlignalTop
BevelOuterbvNoneTabOrder 
DesignSize��   TLabelInstructionsLabelLeftTopWidth�Height'AnchorsakLeftakTopakRight AutoSizeCaption�Instructions for authentication. Please fill in your credentials carefully. Enter all required information, including your session username and session password.XFocusControlPromptEdit1WordWrap	  TLabelPromptLabel1LeftTop8Width�HeightAnchorsakLeftakTopakRight AutoSizeCaption&UsernameX:FocusControlPromptEdit1WordWrap	  TLabelPromptLabel2LeftTopgWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaption&PasswordX:FocusControlPromptEdit2WordWrap	  TPasswordEditPromptEdit1LeftTopJWidth�HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPasswordEditPromptEdit2LeftTopyWidth�HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder   TPanelSavePasswordPanelLeft Top� Width�HeightAlignalTop
BevelOuterbvNoneTabOrder 	TCheckBoxSavePasswordCheckLeftTopWidthHeightCaption   &Ändra lösenord till det härChecked	State	cbCheckedTabOrder    TPanelButtonsPanelLeft Top� Width�Height)AlignalTop
BevelOuterbvNoneTabOrder
DesignSize�)  TButtonPasswordOKButtonLeft� TopWidthPHeightAnchorsakTopakRight CaptionOKModalResultTabOrder   TButtonPasswordCancelButtonLeft� TopWidthPHeightAnchorsakTopakRight CaptionAvbrytModalResultTabOrder  TButtonPasswordHelpButtonLeftHTopWidthPHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick   TPanelSessionRememberPasswordPanelLeft Top� Width�HeightAlignalTop
BevelOuterbvNoneTabOrder 	TCheckBoxSessionRememberPasswordCheckLeftTopWidthHeightCaption.   &Kom ihåg lösenordet för den här sessionenChecked	State	cbCheckedTabOrder     TPanelBannerPanelLeft Top*Width�HeightRAlignalBottom
BevelOuterbvNoneTabOrderVisible
DesignSize�R  TMemo
BannerMemoLeftTopWidth�Height#AnchorsakLeftakTopakRightakBottom Color	clBtnFace	PopupMenuBannerPopupMenuReadOnly	
ScrollBars
ssVerticalTabOrder WantReturnsOnContextPopupBannerMemoContextPopup  	TCheckBoxNeverShowAgainCheckLeftTop7Width� HeightAnchorsakLeftakRightakBottom Caption&   &Visa aldrig det här meddelandet igenTabOrder  TButtonBannerCloseButtonLeft� Top1WidthPHeightAnchorsakRightakBottom Caption	   FortsättModalResultTabOrder  TButtonBannerHelpButtonLeftHTop1WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TActionList
ActionListLeft Top0 	TEditCopyEditCopyActionCategoryBannerCaptionK&opiera
ImageIndex ShortCutC@  TEditSelectAllEditSelectAllActionCategoryBannerCaption&Markera allt
ImageIndexShortCutA@  TActionBannerMonospacedFontActionCategoryBannerCaption   Använd typsnitt &Monospaced	OnExecute!BannerMonospacedFontActionExecute  TActionLabelCopyActionCategoryLabelCaptionK&opiera	OnExecuteLabelCopyActionExecute  TActionLabelOpenLinkAction2CategoryLabelCaption   &Öppna länk	OnExecuteLabelOpenLinkAction2Execute   
TPopupMenuBannerPopupMenuLeft� Top0 	TMenuItemCopyItemActionEditCopyAction  	TMenuItemSelectAllItemActionEditSelectAllAction  	TMenuItemN1Caption-  	TMenuItemAdjustWindowItemActionBannerMonospacedFontAction   
TPopupMenuLabelPopupMenuLeft8TopH 	TMenuItemCopy1ActionLabelCopyAction  	TMenuItemN2Caption-  	TMenuItemOpen1ActionLabelOpenLinkAction2Default	    TPF0TCleanupDialogCleanupDialogLeftdTop� HelpType	htKeywordHelpKeyword
ui_cleanupBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRensa applikationsdataClientHeightCClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnShowFormShow
DesignSize�C 
TextHeight TLabelLabel1LeftTopWidth�HeightlAnchorsakLeftakTopakRight AutoSizeCaption8  Följande lista innehåller all data som det här programmet lagrar på den här datorn. Välj det som du vill ska tas bort.

Om ytterligare instanser av programmet är igång, var god avsluta dem innan nedanstående data tas bort.

Notera att en del av dessa data kommer att återskapas vid nästa uppstart.ShowAccelCharWordWrap	  TButtonOKButtonLeft� Top"WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft=Top"WidthPHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  	TListViewDataListViewLeftTopuWidth�Height� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsCaptionDataWidth�  CaptionPlatsWidth�  ColumnClickDoubleBuffered	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedParentShowHintShowHint	TabOrder 	ViewStylevsReport	OnInfoTipDataListViewInfoTipOnKeyUpDataListViewKeyUpOnMouseDownDataListViewMouseDown  TButtonCheckAllButtonLeftTop"WidthxHeightAnchorsakLeftakBottom CaptionMarkera &allaTabOrderOnClickCheckAllButtonClick  TButton
HelpButtonLeft�Top"WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPF0TConsoleDialogConsoleDialogLeft]Top� HelpType	htKeywordHelpKeyword
ui_consoleBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionKonsolClientHeight�ClientWidth'Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidth�Font.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 	Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�                            (&$�D@=�C@<�C?<�B?<�B>;�A>;�A=:�@=:�@<9�?<9�?;8�>;8�>:7�=:7�=:7�<96�<96�;85�;85�:74�974�963�963�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�.,)�.+)�-+)�-*(�,*(�,)'�+)'�+(&�*(&�*'%�)'%�(&$�(&$�(&$�                            (&$�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�974�963�863�852�752�741�631�630�530�52/�42/�41.�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�.,)�.+)�-+)�,*(�,*(�,)'�+)'�*(&�*(&�)'%�)'%�(&$�(&$�                            (&$�EA>�DA=�D@=�C@<�B?<�B?;�B>;�A>:�@=:�@=:�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�742�741�631�630�520�52/�41/�41.�30.�30-�20-�1/-�1/,�1.,�0.+�/-+�/-*�.,*�.,)�-+)�-+(�,*(�,*'�+)'�+)&�*(&�*(&�)'%�)'%�(&$�                            (&$�EA>�DA>�DA=�C@=�C@<�B?<�B?;�A>;�A>:�@=:�@=9�?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�741�741�631�530�520�52/�41/�31.�30.�20-�2/-�1/,�1.,�0.,�0-+�/-+�/-*�.,*�.,)�-+)�-*(�,*(�,)'�+)'�+)&�*(&�*(&�)'%�(&$�                            (&$�EB>�EA>�DA=�D@=�C@<�C?<�B?<�B>;�A>;�A>:�@=:�@<9�?<9�?;8�>;8�>:7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�.,)�.+)�-+)�-*(�,*(�,)'�+)'�+(&�*(&�*'%�(&$�                            (&$�FB?�EB>�EA>�DA=�D@=�|zw�����usp�B>;�A>;�A=:�@=:�@<9�?<9�>;8�>;8�>:7�=:7�<96�<96�;85�;85�:74�:74�974�963�863�852�752�741�641�630�530�52/�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�.,)�.+)�-+)�-*(�,*(�,)'�+)'�*(&�*(&�(&$�                            (&$�FC?�FB?�EB>�EA>�PMI�����������������QMJ�A>:�@=:�@=:�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�742�741�631�630�520�52/�41/�41.�31.�30-�20-�1/-�1/,�1.,�0.+�/-+�/-*�.,*�.,)�.+)�-+(�,*(�,*'�+)'�+)'�*(&�(&$�                            (&$�GC?�FB?�FB>�EB>�KHE�������������������������A>:�@=:�@=9�?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�742�741�631�630�520�52/�41/�31.�30.�20-�2/-�1/-�1.,�0.,�0.+�/-+�/-*�.,*�.,)�-+)�-*(�,*(�,*'�+)'�+)&�(&$�                            (&$�GC@�FC?�FB?�EB>�EA>�jhd�������������������������YWS�@=:�@<9�?<9�?;8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�752�741�741�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�.,*�.+)�-+)�-*(�,*(�,)'�+)'�(&$�                            (&$�GD@�GC@�FC?�FB?�EB>�EA>�HEA�����������������������������A>;�@<9�?<9�?;8�>;8�>:7�=:7�<96�<96�;85�;85�;85�:74�974�963�863�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�.,)�.+)�-+)�-*(�,*(�,)'�(&$�                            (&$�HD@�GD@�GC@�FC?�FB?�EB>�EA>�DA=�da^�������������������������b`]�@<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�752�741�631�630�520�52/�42/�41.�31.�30-�20-�2/-�1/,�1.,�0.+�/-+�/-*�.,*�.,)�.+)�-+(�,*(�,*(�(&$�                            (&$�HDA�HD@�GC@�GC?�FC?�FB>�EB>�DA>�DA=�EA>�����������������������������EB?�?<8�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�853�852�742�741�631�630�520�52/�41/�31.�30.�30-�2/-�1/-�1/,�0.,�0.+�/-+�/-*�.,*�.,)�-+)�-+(�,*(�(&$�                            (&$�IEA�HDA�HD@�GC@�FC?�FB?�EB>�EA>�DA>�D@=�C@=�XVR�������������������������?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�752�741�741�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-+�/,*�.,*�.,)�-+)�-*(�(&$�                            (&$�IEB�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�[XU���������������������@<9�?<9�?;8�>;8�>:7�=:7�<96�<96�<96�;85�;85�:74�974�963�863�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�.,)�.+)�-+)�(&$�                            (&$�IFB�IEA�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�EB>�����������������������������@=:�@<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�863�852�752�741�631�630�520�52/�42/�41.�31.�30.�20-�2/-�1/,�1.,�0.+�/-+�/-*�/,*�.,)�.+)�(&$�                            (&$�JFB�IEB�IEA�HDA�HD@�GC@�GC?�FC?�FB>�fda�������������������������b_]�A>:�@=:�@=9�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�742�741�631�630�520�52/�41/�41.�30.�30-�2/-�1/-�1/,�0.,�0.+�/-+�/-*�.,*�.,)�(&$�                            (&$�JFC�JFB�IEB�IEA�HDA�HD@�GC@�LIE�����������������������������C@=�B?;�A>;�A>:�@=:�@=9�?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�741�741�631�530�520�52/�41/�31.�30.�20-�2/-�1/,�1.,�0.,�0-+�/-+�/,*�.,*�(&$�                            (&$�JGC�JFB�IFB�IEB�HEA�HDA�vtq�������������������������YVS�C@<�C?<�B?<�B>;�A>;�A>:�@=:�@<9�?<9�?;8�>;8�>:7�=:7�=:7�<96�<96�;85�;85�:74�974�963�963�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�/,*�(&$�                            (&$�KGC�JGC�JFB�IFB�IEB�����������������������������EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�>;8�>;8�>:7�=:7�<96�<96�;85�;85�:74�:74�974�963�863�852�752�741�631�630�530�52/�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�0-+�/-*�(&$�                            (&$�KHD�KGC�JGC�JFB�ZVT���������������������SPL�FB?�EB>�EA>�DA=�D@=�C@<�B?<�B?;�B>;�A>:�@=:�@=:�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�742�741�631�630�520�52/�41/�41.�30.�30-�20-�1/-�1/,�1.,�0.+�/-+�(&$�                            (&$�LHD�KGD�KGC�JFC�MIE�������������ywt�GC@�GC?�FB?�FB>�EA>�DA>�DA=�C@=�C@<�B?<�B?;�A>;�A>:�@=:�@=9�?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�742�741�631�530�520�52/�41/�31.�30.�20-�2/-�1/-�1.,�0.,�0-+�(&$�                            (&$�LHD�KHD�KGC�KGC�JFB�QOK�wtr�NKG�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@=�C?<�B?<�B>;�A>;�A>:�@=:�@<9�?<9�?;8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�0.+�(&$�                            (&$�LIE�LHD�KHD�KGC�JGC�JFB�IFB�IEB�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�>;8�>;8�>:7�=:7�<96�<96�;85�;85�;85�:74�974�963�863�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�2/-�1/,�1.,�(&$�                            (&$�MIE�LIE�LHD�KHD�KGC�JGC�JFB�IEB�IEA�HEA�HD@�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�@=:�@=:�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�752�741�631�630�520�52/�41/�41.�31.�30-�20-�2/-�1/,�(&$�                            (&$�MIE�MIE�LHE�LHD�KGD�KGC�JFC�JFB�IEB�IEA�HDA�HD@�GC@�GC?�FB?�FB>�EB>�DA>�DA=�D@=�C@<�B?<�B?;�A>;�A>:�@=:�@=9�?<9�?<8�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�742�741�631�630�520�52/�41/�31.�30.�20-�2/-�1/-�(&$�                            (&$�NJF�MIE�MIE�LHD�LHD�KGC�KGC�JFC�IFB�IEB�HEA�HDA�HD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@=�C?<�B?<�B?;�A>;�A>:�@=:�@<9�?<9�?;8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�752�741�741�630�530�520�42/�41/�31.�30.�20-�2/-�(&$�                            (&$�NJF�MJF�MIE�MIE�LHD�KHD�KGC�JGC�JFB�IFB�IEB�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�?;8�>;8�>:7�=:7�<96�<96�;85�;85�;85�:74�974�963�863�852�752�741�641�630�530�520�42/�41/�31.�30.�20-�(&$�                            (&$�NJF�NJF�MJF�MIE�LIE�LHD�KHD�KGC�JGC�JFB�IFB�IEA�HEA�HD@�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�@=:�@=:�@<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�752�741�631�630�520�52/�42/�41.�31.�30-�(&$�                            (&$�OKG�NJF�NJF�MIE�MIE�LHE�LHD�KGD�KGC�JGC�JFB�IEB�IEA�HDA�HD@�GC@�GC?�FC?�FB>�EB>�DA>�DA=�D@=�C@<�B?<�B?;�A>;�A>:�@=:�@=9�?<9�?<8�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�853�852�742�741�631�630�520�52/�41/�31.�30.�(&$�                            (&$�OKG�OKG�NJF�NJF�MIE�MIE�LHD�LHD�KGC�KGC�JFC�IFB�IEB�IEA�HDA�HD@�GC@�FC?�FB?�EB>�EA>�DA>�D@=�C@=�C@<�B?<�B?;�A>;�A>:�@=:�@<9�?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�741�741�630�530�520�42/�41/�31.�(&$�                            (&$�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LHD�KHD�KGC�JGC�JFB�IFB�IEB�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�?;8�>;8�>:7�=:7�<96�<96�<96�;85�;85�:74�974�963�863�852�752�741�641�630�530�520�42/�41/�(&$�                            (&$�OKG�OKG�OKG�NJF�NJF�MJF�MIE�LIE�LHD�KHD�KGC�JGC�JFB�IFB�IEA�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�863�852�752�741�631�630�530�52/�42/�(&$�                            (&$�OKG�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LHE�LHD�KGD�KGC�JGC�JFB�IEB�IEA�HDA�HD@�GD@�GC?�FC?�FB>�EB>�EA>�DA=�D@=�C@<�B?<�B?;�B>;�A>:�@=:�@=9�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�742�741�631�630�520�52/�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LHD�LHD�KGD�KGC�JFC�JFB�IEB�IEA�HDA�HD@�GC@�FC?�FB?�FB>�EA>�DA>�DA=�C@=�C@<�B?<�B?;�A>;�A>:�@=:�@=9�?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�741�741�631�530�520�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LHD�KHD�KGC�KGC�JFB�IFB�IEB�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?<�B>;�A>;�A>:�@=:�@<9�?<9�?;8�>;8�>:7�=:7�=:7�<96�<96�;85�;85�:74�974�963�963�852�752�741�641�630�530�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�OKG�OKG�NJF�MJF�MIE�LIE�LHD�KHD�KGC�JGC�JFB�IFB�IEB�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�>;8�>;8�>:7�=:7�<96�<96�;85�;85�:74�:74�974�963�863�852�752�741�631�630�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LHE�LHD�KHD�KGC�JGC�JFB�IEB�IEA�HDA�HD@�GD@�GC?�FC?�FB?�EB>�EA>�DA=�D@=�C@<�B?<�B?;�B>;�A>:�@=:�@=:�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�742�741�631�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LHE�LHD�KGD�KGC�JFC�JFB�IEB�IEA�HDA�HD@�GC@�GC?�FB?�FB>�EB>�DA>�DA=�C@=�C@<�B?<�B?;�A>;�A>:�@=:�@=9�?<9�?<8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�852�742�741�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LHD�KHD�KGC�KGC�JFB�IFB�IEB�HEA�HDA�HD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@=�C?<�B?<�B?;�A>;�A>:�@=:�@<9�?<9�?;8�>;8�>;7�=:7�=:7�<96�<96�;85�;85�:74�:74�963�963�852�752�741�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�NJF�MJF�MIE�LIE�LHD�KHD�KGC�JGC�JFB�IFB�IEB�HEA�HDA�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�A=:�@=:�@<9�?<9�?;8�>;8�>:7�=:7�<96�<96�;85�;85�;85�:74�974�963�863�852�752�(&$�                            (&$�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�OKG�NJF�NJF�MIE�MIE�LIE�LHD�KHD�KGC�JGC�JFB�IEB�IEA�HEA�HD@�GD@�GC@�FC?�FB?�EB>�EA>�DA=�D@=�C@<�C?<�B?;�B>;�A>;�@=:�@=:�?<9�?<9�>;8�>;8�=:7�=:7�<96�<96�;85�;85�:74�:74�964�963�853�852�(&$�                            Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�Ҧ#�                            ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�ӫ%�                            հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�հ'�                            ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�ִ*�                            ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�ع,�                            پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�                            ��0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0���0�                            ��2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �������������������������������������������������      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      ����������������������������������������������������������������(   0   `          �%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              !!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!!                       (&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�###                    (&$�=97�@=:�?<:�?<9�><8�>;8�>:7�=:6�<96�;85�;85�:74�963�963�852�741�641�630�520�420�42/�41/�31.�20-�2/-�1/,�0.+�0-+�/-*�.,)�.+)�-+(�,*(�+)'�+(&�*(&�)'%�)'%�)'%�(&$�(&$�###                    (&$�?<8�D@=�C@<�B?;�A>;�A>:�@=:�?<9�?;8�>;8�=:7�<96�<96�;85�:74�:74�963�853�852�741�631�530�52/�41/�31.�30-�2/-�1/,�1.,�0-+�/-*�.,*�.+)�-+)�,*(�,)'�+)'�*(&�)'%�)'%�(&$�###                    (&$�@<9�DA=�C@=�C?<�B?;�A>;�A=:�@=9�?<9�>;8�>;7�=:7�<96�<96�;85�:74�974�963�852�752�741�630�530�52/�41/�31.�20-�2/-�1/,�0.+�0-+�/-*�.,*�.+)�-*(�,*(�+)'�+)&�*(&�)'%�(&$�###                    (&$�B?;�EA>�DA=�C@<�]ZW�B?;�A>;�@=:�@<9�?<9�>;8�>:7�=:7�<96�;85�;85�:74�964�963�852�752�741�630�520�42/�41.�30.�20-�2/-�1.,�0.+�/-+�/,*�.,)�-+)�-*(�,*(�+)'�*(&�)'%�(&$�###                    (&$�C?<�EB>�DA>�������������ZWT�A>:�@=:�@<9�?<8�>;8�=:7�=:7�<96�;85�;85�:74�963�963�852�741�641�630�520�42/�31.�30.�20-�1/,�1.,�0.+�/-+�/,*�.,)�-+)�,*(�,*'�+)'�)'%�(&$�###                    (&$�C@<�FB?�EB>���������������������DA=�@=:�?<9�?;8�>;8�=:7�<96�<96�;85�:74�:74�963�863�852�741�631�530�52/�41/�31.�30.�2/-�1/,�1.,�0-+�/-*�.,*�.+)�-+)�,*(�,)'�*(&�(&$�###                    (&$�D@=�FC?�FB>�FB?���������������������fca�@=9�?<9�>;8�>;7�=:7�<96�<96�;85�:74�:74�963�852�752�741�631�530�52/�41/�31.�20-�2/-�1/,�0.,�0-+�/-*�.,*�.+)�-+(�,*(�*(&�(&$�###                    (&$�EA=�GC@�FC?�EB>�EA>�XUQ���������������������FB?�?<9�>;8�>:7�=:7�<96�;85�;85�:74�974�963�852�752�741�630�520�42/�41/�30.�20-�2/-�1.,�0.+�/-+�/,*�.,)�-+)�-*(�+)'�(&$�###                    (&$�EA>�GD@�GC?�FB?�EB>�DA>�D@=��~{�����������������olj�?<8�>;8�=:7�=:7�<96�;85�;85�:74�963�963�852�742�641�630�520�42/�41.�30.�20-�1/-�1.,�0.+�/-+�/,*�.,)�-+)�+)'�(&$�###                    (&$�FB>�HDA�GD@�FC?�FB?�EB>�DA=�D@=�OLH�����������������?<9�?;8�>;8�=:7�<96�<96�;85�;85�:74�963�863�852�741�631�530�520�41/�31.�30.�2/-�1/,�1.,�0-+�/-*�.,*�.+)�,*(�(&$�###                    (&$�FB?�HEA�HD@�GC@�FC?�FB>�EA>�KHD���������������������@=9�?<9�>;8�>;8�=:7�<96�<96�;85�:74�:74�963�853�752�741�631�530�52/�41/�31.�30-�2/-�1/,�0.,�0-+�/-*�.,*�-*(�(&$�###                    (&$�GC?�IEB�HEA�HD@�GC@�FC?�zxu�����������������}zx�A>;�@=:�@<9�?<9�>;8�>:7�=:7�<96�<96�;85�:74�974�963�852�752�741�630�520�42/�41/�30.�20-�2/-�1.,�0.+�/-+�/,*�-+(�(&$�###                    (&$�GC@�IFB�IEA�HDA�URO���������������������MJF�B?<�B>;�A>:�@=:�@<9�?<9�>;8�=:7�=:7�<96�;85�;85�:74�964�963�852�742�641�630�520�42/�41.�30.�20-�1/-�1.,�0.+�/-+�.+)�(&$�###                    (&$�HD@�JFB�IFB�yvs�����������������qol�DA=�D@=�C@<�B?<�B>;�A>:�@=:�?<9�?;8�>;8�=:7�=:7�<96�;85�;85�:74�963�863�852�741�631�530�520�41/�31.�30.�2/-�1/,�1.,�0-+�.,)�(&$�###                    (&$�HDA�KGC�JFB�����������������JGC�FB>�EA>�DA=�D@=�C?<�B?;�A>;�A=:�@=:�?<9�>;8�>;8�=:7�<96�<96�;85�:74�:74�963�853�752�741�631�530�52/�41/�31.�30-�2/-�1/,�0.,�/,*�(&$�###                   (&$�IEA�KGC�JGC�fb_�����geb�HD@�GC@�FC?�EB>�EA>�DA=�C@=�C?<�B?;�A>;�@=:�@<9�?<9�>;8�>;7�=:7�<96�<96�;85�:74�974�963�852�752�741�630�520�52/�41/�30.�20-�2/-�1.,�/-*�(&$�###                
(&$�IEB�LHD�KGC�JGC�IFB�IEA�HDA�GD@�GC?�FB?�EB>�EA>�D@=�C@<�B?<�B>;�A>;�@=:�@<9�?<9�>;8�=:7�=:7�<96�;85�;85�:74�964�963�852�742�641�630�520�42/�41.�30.�20-�1/-�0-+�(&$�###                ###(&$�JFB�LHD�KHD�KGC�JFB�IFB�IEA�HDA�GD@�FC?�FB?�EB>�DA>�D@=�C@<�B?<�B>;�A>:�@=:�?<9�?<8�>;8�=:7�=:7�<96�;85�;85�:74�963�863�852�741�631�630�520�41/�31.�30.�20-�0.+�(&$�###                ###(&$�JFB�MIE�LHD�KHD�KGC�JFB�IEB�HEA�HDA�GC@�FC?�FB?�EA>�DA=�D@=�C?<�B?;�A>;�A=:�@=:�?<9�>;8�>;8�=:7�<96�<96�;85�:74�:74�963�853�752�741�631�530�52/�41/�31.�30-�1.,�(&$�###                ###(&$�KGC�MIE�MIE�LHD�KGC�JGC�JFB�IEB�HEA�HD@�GC@�FC?�FB>�EA>�DA=�C@=�C?<�B?;�A>;�@=:�@=9�?<9�>;8�>;7�=:7�<96�<96�;85�:74�974�963�852�752�741�630�520�52/�41/�31.�1/,�(&$�###                ###(&$�KGC�NJF�MIE�LIE�LHD�KGC�JGC�IFB�IEB�HDA�GD@�GC@�FB?�EB>�EA>�D@=�C@<�B?<�B>;�A>;�@=:�@<9�?<9�>;8�>:7�=:7�<96�;85�;85�:74�964�963�852�742�641�630�520�42/�41.�2/-�(&$�###                ###(&$�KHD�NJF�NJF�MIE�LHD�KHD�KGC�JFC�IFB�IEA�HDA�GD@�GC?�FB?�EB>�DA>�D@=�C@<�B?<�B>;�A>:�@=:�?<9�?<8�>;8�=:7�=:7�<96�;85�;85�:74�963�863�852�741�631�630�520�42/�20-�(&$�###                ###(&$�KHD�OKG�NJF�MJF�MIE�LHD�KHD�KGC�JFB�IEB�HEA�HDA�GC@�FC?�FB?�EA>�DA=�D@=�C?<�B?;�A>;�A>:�@=:�?<9�?;8�>;8�=:7�<96�<96�;85�:74�:74�963�853�752�741�631�530�52/�30.�(&$�###                ###(&$�KHD�OKG�OKG�NJF�MIE�MIE�LHD�KGD�JGC�JFB�IEB�HEA�HD@�GC@�FC?�FB>�EA>�DA=�C@=�C?<�B?;�A>;�@=:�@=9�?<9�>;8�>;7�=:7�<96�<96�;85�:74�974�963�852�752�741�630�530�41.�(&$�###                ###(&$�KHD�OKG�OKG�OKG�NJF�MIE�LIE�LHD�KGC�JGC�IFB�IEB�HDA�GD@�GC@�FB?�EB>�EA>�D@=�C@<�B?<�B?;�A>;�@=:�@<9�?<9�>;8�>:7�=:7�<96�;85�;85�:74�964�963�852�742�741�630�41/�(&$�###                ###(&$�KHD�OKG�OKG�OKG�NJF�NJF�MIE�LHE�KHD�KGC�JFC�IFB�IEA�HDA�GD@�GC?�FB?�EB>�DA>�D@=�C@<�B?<�B>;�A>:�@=:�@<9�?<8�>;8�=:7�=:7�<96�;85�;85�:74�963�863�852�741�641�42/�(&$�###                ###(&$�KHD�OKG�OKG�OKG�OKG�NJF�MJF�MIE�LHD�KHD�KGC�JFB�IEB�HEA�HDA�GC@�FC?�FB?�EA>�DA=�D@=�C@<�B?;�A>;�A>:�@=:�?<9�?;8�>;8�=:7�<96�<96�;85�:74�:74�963�853�852�741�420�(&$�###                ###(&$�KHD�OKG�OKG�OKG�OKG�OKG�NJF�MIE�MIE�LHD�KGD�JGC�JFB�IEB�HEA�HD@�GC@�FC?�FB>�EA>�DA=�C@=�C?<�B?;�A>;�A=:�@=9�?<9�>;8�>;7�=:7�<96�<96�;85�:74�974�963�852�752�520�(&$�###                ###(&$�KHD�OKG�OKG�OKG�OKG�OKG�OKG�NJF�MIE�LIE�LHD�KGC�JGC�IFB�IEB�HDA�HD@�GC@�FB?�EB>�EA>�DA=�C@<�B?<�B?;�A>;�@=:�@<9�?<9�>;8�>:7�=:7�<96�;85�;85�:74�964�963�852�520�(&$�
                ###(&$�KHD�OKG�OKG�OKG�OKG�OKG�OKG�NJF�NJF�MIE�LHE�KHD�KGC�JFC�IFB�IEA�HDA�GD@�GC?�FB?�EB>�DA>�D@=�C@<�B?<�B>;�A>:�@=:�@<9�?<8�>;8�=:7�=:7�<96�;85�;85�:74�963�963�630�(&$�                    ###ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�ҧ#�                    ###ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�ԭ&�                       ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�ִ)�                        غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�غ,�                        ��/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/�                        ��2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ������  ������  ������  ������  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      ������  ������  ������  ������  ������  ������  (   (   P          @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�                (&$�D@=�C@<�B?;�A>;�@=:�@<9�?<8�>;8�=:7�<96�;85�;85�:74�963�853�752�741�630�520�41/�31.�20-�2/-�1.,�0.+�/-*�.,*�.+)�-*(�,*'�+)'�*(&�)'%�(&$�(&$�                (&$�DA=�D@=�C?<�B?;�A>;�@=:�?<9�?;8�>;7�=:7�<96�;85�;85�:74�963�852�742�641�530�52/�41/�30.�20-�1/-�1.,�0-+�/-*�.,)�-+)�,*(�,)'�+)&�*(&�)'%�(&$�                (&$�EB>�DA=�JGD�����jgd�A>:�@=:�?<9�>;8�>:7�=:7�<96�;85�:74�974�963�852�741�631�530�52/�41/�30.�20-�1/,�0.,�0-+�/,*�.,)�-+)�,*(�,)'�+(&�*(&�(&$�                (&$�FB?�EA>�pnk�������������JFC�@=9�?<9�>;8�=:7�=:7�<96�;85�:74�964�963�852�741�630�520�42/�31.�30.�2/-�1/,�0.+�/-+�/,*�.,)�-+(�,*(�+)'�*(&�(&$�                (&$�FC?�FB>�EA>�����������������xvt�@<9�?<9�>;8�=:7�<96�<96�;85�:74�963�853�752�741�630�520�42/�31.�30-�2/-�1.,�0.+�/-*�.,*�.+)�-*(�,*(�+)'�(&$�                (&$�GC@�FC?�EB>�DA>�YVS�����������������OKH�?;8�>;8�=:7�<96�;85�;85�:74�963�852�752�641�630�520�41/�31.�20-�1/-�1.,�0-+�/-*�.,*�-+)�-*(�,)'�(&$�                (&$�HD@�GC@�FB?�EB>�DA=�C@=����������������omk�>;8�>;7�=:7�<96�;85�:74�:74�963�852�742�631�530�52/�41/�30.�20-�1/,�1.,�0-+�/-*�.,)�-+)�,*(�(&$�                (&$�HEA�GD@�GC?�FB?�EA>�DA=�JGC�����������������?<9�>;8�>:7�=:7�<96�;85�:74�974�963�852�741�631�530�42/�41.�30.�2/-�1/,�0.+�/-+�/,*�.,)�-+)�(&$�                (&$�IEB�HDA�GD@�FC?�FB>�yvt�����������������B>;�@=9�?<9�>;8�=:7�<96�<96�;85�:74�963�863�852�741�630�520�42/�31.�30-�2/-�1/,�0.+�/-+�.,*�.+)�(&$�                (&$�IFB�IEA�HDA�URO�����������������XVR�B?;�A>;�@=:�@<9�?<8�>;8�=:7�<96�;85�;85�:74�963�853�752�741�630�520�41/�31.�20-�2/-�1.,�0.+�/-*�.,*�(&$�                (&$�JFC�IFB�`^Z�����������������DA=�D@=�C?<�B?;�A>;�@=:�?<9�?;8�>;7�=:7�<96�;85�;85�:74�963�852�742�641�630�52/�41/�30.�20-�1/-�1.,�0-+�/-*�(&$�                (&$�KGC�JFB�c_]���������TPL�FB?�EB>�DA=�C@=�B?<�B>;�A>:�@=:�?<9�>;8�>:7�=:7�<96�;85�:74�974�963�852�741�631�530�52/�41/�30.�20-�1/,�0.,�0-+�(&$�                (&$�KHD�KGC�JFB�IEB�HDA�GD@�FC?�FB?�EA>�DA=�C@<�B?<�B>;�A>:�@=9�?<9�>;8�=:7�=:7�<96�;85�:74�964�963�852�741�631�520�42/�31.�30.�2/-�1/,�0.+�(&$�                (&$�LHD�KGD�JGC�JFB�IEA�HDA�GC@�FC?�FB>�EA>�D@=�C@<�B?;�A>;�@=:�@<9�?<9�>;8�=:7�<96�<96�;85�:74�963�853�752�741�630�520�42/�31.�30-�2/-�1.,�(&$�                (&$�MIE�LHD�KGC�JGC�IFB�IEA�HDA�GC@�FC?�EB>�DA>�D@=�C?<�B?;�A>;�@=:�@<9�?;8�>;8�=:7�<96�;85�;85�:74�963�852�752�741�630�520�41/�31.�20-�1/-�(&$�                (&$�MIE�MIE�LHD�KGC�JFC�IEB�HEA�HD@�GC@�FB?�EB>�DA=�C@=�C?<�B?;�A>:�@=:�?<9�>;8�>;7�=:7�<96�;85�:74�:74�963�852�742�631�530�52/�41/�30.�20-�(&$�                (&$�NJF�MIE�LIE�KHD�KGC�JFB�IEB�HEA�GD@�GC?�FB?�EA>�DA=�C@<�B?<�B>;�A>:�@=:�?<9�>;8�>:7�=:7�<96�;85�:74�974�963�852�741�631�530�42/�41.�30.�(&$�                (&$�OKG�NJF�MIE�LHD�KHD�KGC�JFB�IEB�HDA�GD@�FC?�FB>�EA>�D@=�C@<�B?<�A>;�A=:�@=9�?<9�>;8�=:7�<96�<96�;85�:74�963�863�852�741�630�520�42/�31.�(&$�                (&$�OKG�NJF�NJF�MIE�LHD�KGD�JGC�IFB�IEA�HDA�GC@�FC?�EB>�EA>�D@=�C@<�B?;�A>;�@=:�@<9�?<8�>;8�=:7�<96�;85�;85�:74�963�853�752�741�630�520�41/�(&$�                (&$�OKG�OKG�NJF�MJF�MIE�LHD�KGC�JFC�IFB�HEA�HD@�GC@�FB?�EB>�DA=�D@=�C?<�B?;�A>;�@=:�?<9�?;8�>;7�=:7�<96�;85�;85�:74�963�852�742�641�630�52/�(&$�                (&$�OKG�OKG�OKG�NJF�MIE�LIE�LHD�KGC�JFB�IEB�HEA�HD@�GC?�FB?�EB>�DA=�C@=�C?<�B>;�A>:�@=:�?<9�>;8�>:7�=:7�<96�;85�:74�974�963�852�741�631�530�(&$�                (&$�OKG�OKG�OKG�OKG�NJF�MIE�LHE�KHD�KGC�JFB�IEB�HDA�GD@�FC?�FB?�EA>�DA=�C@<�B?<�B>;�A>:�@=9�?<9�>;8�=:7�=:7�<96�;85�:74�964�963�852�741�631�(&$�                (&$�OKG�OKG�OKG�OKG�OKG�NJF�MIE�LHD�KGD�JGC�JFB�IEA�HDA�GC@�FC?�FB>�EA>�D@=�C@<�B?;�A>;�@=:�@<9�?<9�>;8�=:7�<96�<96�;85�:74�963�863�752�741�(&$�                (&$�OKG�OKG�OKG�OKG�OKG�NJF�MJF�MIE�LHD�KGC�JGC�IFB�IEA�HDA�GC@�FC?�EB>�DA>�D@=�C?<�B?;�A>;�@=:�@<9�?;8�>;8�=:7�<96�;85�;85�:74�963�852�752�(&$�                (&$�OKG�OKG�OKG�OKG�OKG�OKG�NJF�MIE�MIE�LHD�KGC�JFC�IEB�HEA�HD@�GC@�FB?�EB>�DA=�D@=�C?<�B?;�A>:�@=:�?<9�>;8�>;7�=:7�<96�;85�:74�:74�963�852�(&$�                Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�Ҩ$�                կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�կ'�                ׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�                پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�پ.�                ��2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2���2�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����   �����   �����   �����   �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �����   �����   �����   �����   �����   (       @          �                                                                                                                                                                                                                                                                                                                                                                                                                      (&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�        (&$�D@=�C?<�B>;�A=:�@<9�?;8�>;7�=:7�<96�;85�:74�963�852�741�630�52/�41/�30.�2/-�1.,�0-+�/,*�.,)�-*(�,*'�+)&�*(&�)'%�(&$�        (&$�DA=�C@=�B?<�A>;�@=:�?<9�>;8�=:7�<96�;85�;85�974�963�752�741�530�52/�31.�30-�1/-�1.,�/-+�/,*�.+)�-*(�,)'�+(&�*'%�(&$�        (&$�EB>�DA=���������MJG�@=:�?<9�>;8�=:7�<96�;85�:74�964�853�752�631�530�42/�31.�20-�1/,�0.+�/-+�.,*�-+)�,*(�+)'�*(&�(&$�        (&$�FB?�EA>�mjh���������}{y�@=9�?<9�>;8�=:7�<96�;85�:74�963�852�741�630�520�41/�30.�20-�1/,�0.+�/-*�.,)�-+)�,*(�+)'�(&$�        (&$�GC?�FB?�EA>�HDA�������������D@=�?;8�>;7�=:7�<96�;85�:74�963�852�741�630�52/�41/�30.�2/-�1.,�0-+�/,*�.,)�-+(�,*'�(&$�        (&$�GD@�FC?�EB>�DA>�������������FC@�?<9�>;8�=:7�<96�;85�;85�974�963�752�741�530�52/�31.�30-�1/-�1.,�/-+�/,*�.+)�-*(�(&$�        (&$�HDA�GD@�_]Y�������������C@<�A>;�@=:�?<9�>;8�=:7�<96�;85�:74�964�853�752�631�530�42/�31.�20-�1/,�0.+�/-+�.,*�-+)�(&$�        (&$�IEB�HDA���������ZVT�DA=�C@<�B?;�A>:�@=:�?<9�>;8�=:7�<96�;85�:74�963�852�741�631�520�41/�30.�20-�1/,�0.+�/-*�.,)�(&$�        (&$�JFB�IEA�QMJ�GC@�FB?�EA>�D@=�C?<�B>;�A>:�@<9�?<8�>;7�=:7�<96�;85�:74�963�852�741�630�520�41/�30.�2/-�1.,�0-+�/-*�(&$�        (&$�JGC�IFB�HEA�GD@�FC?�EB>�DA>�D@=�B?<�B>;�@=:�@<9�>;8�>:7�<96�<96�;85�:74�963�852�741�630�52/�41.�30-�2/-�1.,�0-+�(&$�        (&$�KGD�JFC�IEB�HDA�GD@�FC?�EB>�DA=�C@<�B?;�A>;�@=:�?<9�>;8�=:7�<96�;85�:74�964�863�752�641�530�42/�31.�20-�1/,�0.,�(&$�        (&$�LHD�KGC�JFB�IEB�HDA�GC@�FB?�EA>�DA=�C@<�B?;�A>:�@=:�?<9�>;8�=:7�<96�;85�:74�963�852�741�631�520�41/�31.�20-�1/,�(&$�        (&$�MIE�LHD�KGC�JFB�IEA�HD@�GC@�FB?�EA>�D@=�C?<�B>;�A>:�@<9�?<8�>;7�=:7�<96�;85�:74�963�852�741�630�520�41/�30.�2/-�(&$�        (&$�MJF�LIE�KHD�JGC�IFB�HEA�HD@�FC?�FB>�DA>�D@=�B?<�B>;�@=:�@<9�>;8�>:7�<96�<96�;85�:74�963�852�741�630�52/�41.�30-�(&$�        (&$�NJF�MIE�LHE�KGD�JGC�IEB�HEA�GD@�FC?�EB>�DA=�C@<�B?<�A>;�@=:�?<9�>;8�=:7�<96�;85�:74�964�863�752�641�530�42/�31.�(&$�        (&$�OKG�NJF�MIE�LHD�KGC�JFB�IEB�HDA�GC@�FB?�EB>�DA=�C@<�B?;�A>;�@=:�?<9�>;8�=:7�<96�;85�:74�963�852�742�631�520�41/�(&$�        (&$�OKG�OKG�NJF�MIE�LHD�KGC�JFB�IEA�HDA�GC@�FB?�EA>�D@=�C?<�B?;�A>:�@=9�?<8�>;8�=:7�<96�;85�:74�963�852�741�630�520�(&$�        (&$�OKG�OKG�NJF�MJF�LIE�KHD�JGC�IFB�HEA�HD@�FC?�FB>�EA>�D@=�C?<�B>;�A=:�@<9�?;8�>:7�=:7�<96�;85�:74�963�852�741�630�(&$�        (&$�OKG�OKG�OKG�NJF�MIE�LHE�KGD�JGC�IEB�HEA�GD@�FC?�EB>�DA=�C@<�B?<�A>;�@=:�?<9�>;8�=:7�<96�;85�:74�974�863�752�641�(&$�        (&$�OKG�OKG�OKG�OKG�NJF�MIE�LHD�KGC�JFB�IEB�HDA�GC@�FB?�EB>�DA=�C@<�B?;�A>;�@=:�?<9�>;8�=:7�<96�;85�:74�963�853�742�(&$�        (&$�OKG�OKG�OKG�OKG�OKG�NJF�MIE�LHD�KGC�JFB�IEA�HDA�GC@�FB?�EA>�D@=�C?<�B?;�A>:�@=9�?<8�>;8�=:7�<96�;85�:74�963�852�(&$�        ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�ө$�        ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�ֲ)�        ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�ټ-�        ��1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1�                                                                                                                                                                                                                                                                                                                                                                                                    �������������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ������������(      0          `	                                                                                                                                                                                                                  (&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�D@=�B?<�A>;�@=9�?;8�=:7�<96�;85�974�853�741�630�42/�30.�2/-�0.,�/-*�.,)�,*(�+)'�*(&�)'%�'%#�(&$�EA>�D@=�ROM�A>:�@<9�>;8�=:7�<96�;85�964�852�741�530�41/�30.�1/-�0.+�/-*�.+)�,*(�+)'�*(&�'%#�(&$�FB?�EA>���������YWS�?<9�>;8�=:7�<96�:74�963�852�641�520�41/�30-�1/,�0.+�/,*�-+)�,*(�+)&�'%#�(&$�GC@�FB?�\YW�������������@=:�>;8�=:7�;85�:74�963�752�631�520�41.�20-�1/,�0-+�.,*�-+)�,*'�'%#�(&$�HDA�GC@�FB>�DA=�������������C@=�>;7�<96�;85�:74�963�752�630�52/�31.�20-�1.,�/-+�.,)�-+(�'%#�(&$�IEB�HDA�GC?�NKG�������������A>;�?<8�=:7�<96�;85�:74�863�741�630�42/�31.�2/-�1.,�/-*�.,)�'%#�(&$�JGC�IEB�|zw���������tqn�B?<�A>;�@=9�>;8�=:7�<96�;85�974�852�741�530�42/�30.�2/-�0.+�/-*�'%$�(&$�KHD�JFB���������LIE�EA>�D@=�B?;�A>:�@<9�>;8�=:7�<96�;85�963�852�741�530�41/�30.�1/,�0.+�'&$�(&$�LIE�KGC�JFB�HEA�GD@�FB?�EA>�C@<�B?;�A=:�?<9�>;8�=:7�<96�:74�963�852�641�520�41/�20-�1/,�(&$�(&$�MJF�LHD�KGC�IFB�HEA�GC@�FB?�DA=�C@<�B>;�@=:�?<9�>;8�<96�;85�:74�963�752�631�520�31.�20-�(&$�(&$�NJF�MIE�LHD�KGC�IFB�HDA�GC@�EB>�DA=�C?<�B>;�@=:�?<9�>:7�<96�;85�:74�963�742�630�52/�31.�(&$�(&$�OKG�NJF�MIE�LHD�JGC�IEB�HDA�FC?�EB>�D@=�C?<�A>;�@=:�?;8�=:7�<96�;85�:74�853�741�630�42/�(&$�(&$�OKG�OKG�NJF�MIE�KHD�JFC�IEB�HD@�FC?�EA>�D@=�B?<�A>;�@<9�>;8�=:7�<96�;85�964�852�741�530�(&$�(&$�OKG�OKG�OKG�NJF�MIE�KGD�JFB�IEA�GD@�FB?�EA>�C@=�B?;�A>:�@<9�>;8�=:7�<96�:74�963�852�741�(&$�(&$�OKG�OKG�OKG�OKG�MJF�LHE�KGC�JFB�HEA�GC@�FB?�DA>�C@<�B?;�A=:�?<9�>;8�=:7�;85�:74�963�852�(&$�(&$�OKG�OKG�OKG�OKG�OKG�MIE�LHD�KGC�IFB�HDA�GC@�FB>�DA=�C@<�B>;�@=:�?<9�>;7�<96�;85�:74�963�(&$�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1�                                                                                                                                                                                                ��� ���                                                                                 ��� ��� (      (          �                                                                                                                                                                                  (&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�D@=�B?;�QNK�?<9�>:7�<96�:74�963�742�630�41/�30-�1.,�/-+�.,)�,*(�+(&�)'%�(&$�(&$�EA>�C@=���������XTR�=:7�<96�:74�863�741�530�41.�20-�1.,�/-*�-+)�,*'�*(&�(&$�(&$�FC?�EA>�XVR�������������>;8�;85�:74�852�641�520�31.�2/-�0.+�/,*�-+)�,)'�(&$�(&$�GD@�FB?�DA=�C?<�������������<96�;85�964�852�631�52/�30.�1/,�0-+�.,*�-*(�(&$�(&$�IEA�GC@�EB>�TPN�������������>:7�<96�:74�963�752�630�41/�30-�1/,�/-+�.,)�(&$�(&$�JFB�HDA�������������b`]�@=:�?<8�=:7�<96�:74�963�741�530�41/�20-�1.,�/-*�(&$�(&$�KGC�IFB���������FB?�C@<�B>;�@=9�>;8�=:7�;85�:74�852�741�520�31.�2/-�0.+�(&$�(&$�LHD�KGC�IEB�GD@�FB?�DA=�C?<�A>;�@<9�>;8�<96�;85�964�852�631�52/�30.�1/-�(&$�(&$�MIE�LHD�JFC�IEA�GC@�EB>�D@=�B?<�A>:�?<9�>:7�<96�;85�963�752�630�42/�30-�(&$�(&$�OKG�MIE�KHD�JFB�HDA�GC?�EB>�D@=�B?;�@=:�?<8�=:7�<96�:74�963�741�530�41/�(&$�(&$�OKG�NJF�MIE�KGC�IFB�HDA�FC?�EA>�C@<�B>;�@=:�>;8�=:7�;85�:74�852�741�520�(&$�(&$�OKG�OKG�NJF�LHD�KGC�IEB�HD@�FB?�DA=�C?<�A>;�@<9�>;8�<96�;85�964�852�631�(&$�(&$�OKG�OKG�OKG�MIE�LHD�JGC�IEA�GC@�FB>�DA=�B?<�A>:�?<9�>:7�<96�;85�963�752�(&$�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�Ӫ%�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+�׷+���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1���1�                                                                                ��� ���                                                                     ��� (                 @                                                                                  (&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�(&$�D@=�D@=�@<9�>:7�<96�:74�852�630�41.�2/-�0-+�.+)�,)'�*(&�(&$�(&$�EB>���������KHE�=:7�;85�963�742�520�31.�1/,�/-*�-+)�+)'�(&$�(&$�GC?�ifd���������|z�=:7�;85�963�741�52/�30.�1.,�/,*�-*(�(&$�(&$�HDA�FC?�GD@�������������<96�:74�853�631�42/�20-�0.+�.,*�(&$�(&$�JFB�HD@�MIF�������������>;7�<96�:74�852�630�41/�2/-�0-+�(&$�(&$�KGD�zwu���������sqn�A>;�?<9�=:7�;85�964�752�530�31.�1/,�(&$�(&$�MIE���������MIE�EA>�C?<�A>:�?<8�=:7�;85�963�741�520�30.�(&$�(&$�NJF�LHD�JFC�HDA�FC?�DA=�B?;�@=:�>;8�<96�:74�863�641�42/�(&$�(&$�OKG�NJF�LHD�JFB�HD@�FB?�D@=�B>;�@<9�>;7�<96�:74�852�630�(&$�(&$�OKG�OKG�MIE�KGD�IEB�GD@�EB>�C@<�A>;�?<9�=:7�;85�964�752�(&$�(&$�OKG�OKG�OKG�MIE�KGC�IEA�GC@�EA>�C?<�A>:�?<8�=:7�;85�963�(&$�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&�Ԯ&���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/���/�                                                                ��                                                          ��  OnCloseQueryFormCloseQueryOnShowFormShow
DesignSize'� 
TextHeight TBevelBevel1Left Top Width'HeightPAlignalTopShapebsBottomLine  TLabelLabel1Left3TopWidthXHeightCaptionAnge &kommando:FocusControlCommandEdit  TLabelLabel2Left3Top8Width]HeightCaptionAktuell katalog:ShowAccelChar  TLabelLabel4Left3Top"Width�HeightAnchorsakLeftakTopakRight AutoSizeCaptionP   Varning: Kör inga kommandon som kräver användardata eller dataöverföringar.ShowAccelChar  
TPathLabelDirectoryLabelLeft� Top8Width*HeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TImageImageLeftTopWidth Height AutoSize	  TMemo
OutputMemoLeft TopPWidth'Height9TabStopAlignalClientColor	clBtnFace	PopupMenu	PopupMenuReadOnly	
ScrollBarsssBothTabOrderWantReturnsOnContextPopupOutputMemoContextPopup  TButton	CancelBtnLeft�TopWidthPHeightAnchorsakTopakRight Cancel	Caption   StängModalResultTabOrder  THistoryComboBoxCommandEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength TabOrder OnChangeCommandEditChange  TButtonExecuteButtonLeftyTopWidthPHeightAnchorsakTopakRight Caption   K&örDefault	TabOrderOnClickExecuteButtonClick  TButton
HelpButtonLeft�Top*WidthPHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TPngImageListImages	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:43+01:00" xmp:MetadataDate="2022-09-01T11:00:43+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9e4a76d0-ec4c-a349-8e28-329bad9961d7" xmpMM:DocumentID="adobe:docid:photoshop:d3f5036e-852f-5349-b6a9-2cdc138995b9" xmpMM:OriginalDocumentID="xmp.did:53c73639-e58b-b149-ae33-49bc5bbe7e24"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:53c73639-e58b-b149-ae33-49bc5bbe7e24" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9e4a76d0-ec4c-a349-8e28-329bad9961d7" stEvt:when="2022-09-01T11:00:43+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>F!�*   �IDATx�c���?��Y��3`��@A����#8 H/#̀��X�9�3���|���'.C�����}���` ��l(�����J��]4��h �8Q��J(f��P�t���JK:'!1��̴$V�����0m�\�14����b�(�� � z���J�xC    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:46+01:00" xmp:MetadataDate="2022-09-01T11:00:46+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a1cb064b-38bb-d143-aca5-917a4f08a7cc" xmpMM:DocumentID="adobe:docid:photoshop:37c98265-f6fc-1b48-998e-ab64cb46ee56" xmpMM:OriginalDocumentID="xmp.did:7460783c-7362-1449-9e0a-d4169f0168f5"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7460783c-7362-1449-9e0a-d4169f0168f5" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a1cb064b-38bb-d143-aca5-917a4f08a7cc" stEvt:when="2022-09-01T11:00:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>b%��  �IDATx�c���?%�d��Y��2%3-�n �C�f��,{��a�ӏ�?�d`��Y������	���g��������������?�����=I�pA��\yΰhH�?C��8�w���#������,��0�R��~C����۟2Ԝ{�p��Ws�E�
� ��������5�����,D�;*�7���s��>00M��f� �C�?3~�l�g%������n�-p�M0�ap�<�{̰��{K	�<����u�m��ی���|������� ���;�?� �Ƞ���p��vf&�/��2���5���}����3�z������!PI��蒊O���(�ɂ?�J�e&J  ���mG�&    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:48+01:00" xmp:MetadataDate="2022-09-01T11:00:48+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:dfee8aa3-ad36-f244-9f21-d3e2e6e2eca3" xmpMM:DocumentID="adobe:docid:photoshop:2600ec29-7b04-494d-919e-8e57935905cc" xmpMM:OriginalDocumentID="xmp.did:d4ca593b-0a91-0a4d-9f68-949bca3e41e4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d4ca593b-0a91-0a4d-9f68-949bca3e41e4" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:dfee8aa3-ad36-f244-9f21-d3e2e6e2eca3" stEvt:when="2022-09-01T11:00:48+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�'ߌ  �IDATx�c���?%�Q��-�M�`��Ȩ��
���fdTQ���������$%0̜5����{��-���Q@V����0���!;�����K(��|��� P`"+���à���p�����\��#���a�����0�ڷ�����v���'��ʪ:�Z���E�pE��a��q �1m2���Μ9����g�uuu�ё(!lc�����C(r�g�b���G ����Cb|,Cn~\���̭l��Y3�1L�>����3߿C +� �7�?�9�`ja�6 ����Ҳ�(!󯾞.�`&���2���a���,�]]��@''��3�;wÅ��F )%�UP�ٙ�'O�0�����0�ܼ 6��� SE�����    IEND�B`�  LeftHTop�   
TPopupMenu	PopupMenuImagesImagesLeft�Top�  	TMenuItemCopyItemActionEditCopy  	TMenuItemSelectAllItemActionEditSelectAll  	TMenuItemN1Caption-  	TMenuItemAdjustWindowItemActionAdjustWindow   TActionList
ActionListImagesImages	OnExecuteActionListExecuteOnUpdateActionListUpdateLeftHTop�  	TEditCopyEditCopyCaptionK&opiera
ImageIndex ShortCutC@  TEditSelectAllEditSelectAllCaption&Markera allt
ImageIndexShortCutA@  TActionAdjustWindowCaption   Anpassa &fönster
ImageIndexShortCutJ@   TPngImageList	Images120HeightWidth	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:43+01:00" xmp:MetadataDate="2022-09-01T11:00:43+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0d3bd438-11f1-7c4d-9bd7-9f4d1f44ec66" xmpMM:DocumentID="adobe:docid:photoshop:f88caac6-6121-fe41-b67a-0914eaa6a23c" xmpMM:OriginalDocumentID="xmp.did:15f53f04-50a4-0841-b549-c1916a4208ba"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:15f53f04-50a4-0841-b549-c1916a4208ba" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0d3bd438-11f1-7c4d-9bd7-9f4d1f44ec66" stEvt:when="2022-09-01T11:00:43+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>e�.   �IDATx�c���?��Y��3������G �Y�0Sc�*�31˗��x2�h}�=���C�PA���?Y�ɬ�ݵ@�v!6גd ]]��$)�c��$E��MRYiIG�v!1I*3-��"/����HD^f 6I�ddę�͜Kt�"��QR�B�H�4(  M ��*    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:46+01:00" xmp:MetadataDate="2022-09-01T11:00:46+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6e475de9-188e-1b46-9896-52eae0273cd8" xmpMM:DocumentID="adobe:docid:photoshop:08154e42-e852-384b-bd56-9e4e94073a78" xmpMM:OriginalDocumentID="xmp.did:81e9d631-92e3-a34b-b0e0-e410f6c9dc99"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:81e9d631-92e3-a34b-b0e0-e410f6c9dc99" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6e475de9-188e-1b46-9896-52eae0273cd8" stEvt:when="2022-09-01T11:00:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Kh�  �IDATxڵ��/�Aǿ�V�J[-UI�Jh�*v�B�"A,�p�!�����Op$ĕd����-ًD��X�R�mV���o��v~�.q2�z��33���|g�g8��N����tZ��}�#�,^#�����?�0��D�<4R1*2��O��a��g�<�% &Y���6����b��q$����?*�[�a��ܘ�{h`�^�A�o�v��7��\��d�{6`��܅q��C��8q9W0���c�ҠȄ�ِZQ��İ�	`�Ī��m�*4
�#;p�V7���=yTʰ��hv�0�㠁"�C�65������g픂��L,���[�m�߅i�\}	�ret�*E�#��\�K+�B���X�j����E1_x���9���$�
����L*l�+�]�G�2��]�8=S�#�z{9���-F6ϚZ��,	$D��|E�o3A�!b������ݴM4ߩ0�Q˹�=3T�ç|yj}�jo|-i��t�?^��:�xI    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
h  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:49+01:00" xmp:MetadataDate="2022-09-01T11:00:49+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0b372f15-4296-ff41-bc3c-129cbae619d8" xmpMM:DocumentID="adobe:docid:photoshop:7d25028b-f463-f843-87fa-9e90ff8f8ca6" xmpMM:OriginalDocumentID="xmp.did:980b368d-d655-6d45-ba5f-8ccdda364327"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:980b368d-d655-6d45-ba5f-8ccdda364327" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0b372f15-4296-ff41-bc3c-129cbae619d8" stEvt:when="2022-09-01T11:00:49+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Y�4  KIDATx�c���?5����T5�Q{�u����2uTQ��������(\��P��ř�`رs\��? ����ç�QDH��� +#�0{�T�|RJ:�����Y���'��`I$��]���
6LNVl��G�S���7��/_>CTRQ��
�֪�7W�0ھc'CCS��|��b���*X����!/7��������p:|`/�0k{�pk��ahm�d����߿}�������*99Ygw��6���%�Ξ:�p�����R����2���b`jZC~N;;;֤`ic6���CX� ô���aժ�SRS
r�qham6���8ljieX�z�@YyE9i�ƆZy99g�wA�t��A�Fs+���p�4ý��

��ܽ����/��2r��dR\����ց�0��Y����z���6��߿�-���7�@iY9����@h���b��pG��֭��jk��#|�����RҲA�l���ưh�\yyy�a��$<*�"l �l����m��t���|��4f���[�H�	���6n"\�P�Ħ�� ���E��    IEND�B`�  Left�Top�   TPngImageList	Images144HeightWidth	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:44+01:00" xmp:MetadataDate="2022-09-01T11:00:44+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e21335c1-f1bb-a24b-9cca-c2be37f8c391" xmpMM:DocumentID="adobe:docid:photoshop:dc254fa2-c914-f74d-bd30-90b824bc6bba" xmpMM:OriginalDocumentID="xmp.did:9cdc2fa1-ceab-004d-b67f-53c9282ab6da"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:9cdc2fa1-ceab-004d-b67f-53c9282ab6da" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e21335c1-f1bb-a24b-9cca-c2be37f8c391" stEvt:when="2022-09-01T11:00:44+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���R   �IDATx�c���?��Y��3��
�ӓ�0� @f3�,HI�ũp���,,,_~���I�%$Y�����}��,!����W�I���A� �����dV�� ���0R��|D���x F^!����O=���R�
�}��W�Ғ���R�JfZ+�|�M=�F�- %��X@����##�<�0m�\�s;Y��`���m:�,  u"i�p>.    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:47+01:00" xmp:MetadataDate="2022-09-01T11:00:47+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8a0ab898-272e-4442-93b1-44f6837fb2be" xmpMM:DocumentID="adobe:docid:photoshop:bfe1f4b8-13f6-2740-a13d-1fcf34f5a993" xmpMM:OriginalDocumentID="xmp.did:d8dc3fe3-1bd0-fb4d-bdaa-bd4f25d9aa67"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d8dc3fe3-1bd0-fb4d-bdaa-bd4f25d9aa67" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8a0ab898-272e-4442-93b1-44f6837fb2be" stEvt:when="2022-09-01T11:00:47+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>?wn$  tIDATx�͕]H�QƟwn�u��9�V��i�
*��(04�o�݅PAw��J��*��
#!���u#	����b}l6��t_�طo�s�^&��N�ag{~�<��	�,��%0��U���w
�&�*N���@z�R9��+k4huh���	��q�A<S Vd�L��Q"�E�	g[�C�0��w��F�|~�n��ͨ�';μ�!��!��A�р:ڵ'��g�p�%���� ̚����}O�`o�������Xp	�2��K�V�Ei����t�.��j�/�T��3W��m��RT�x���X
��I��%J攞��"@}�i��e ���$��7�hKy�]�6�� ���y<��)6��F�fQ��hJI�H�J�c�x`f^�I"�Zp�Tǽ~���_��ho�:��7��]�rq�Z���0PDK�����A.�J5`���Qv��M<<ֺj��۟x5W���=����[��{��{3�5
�d ��%/����X�~��O!{��Ŀkv�h,��dvM���N4K�,f�����rVi$�c�F���;10�++��ء�D�����qz�I��Q�V��M� �n�������)�W�6R�����R լ?&����    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:50+01:00" xmp:MetadataDate="2022-09-01T11:00:50+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:7af6382a-5db8-f840-b3e3-149686d7e425" xmpMM:DocumentID="adobe:docid:photoshop:061ca7f5-0366-db43-9c6b-6e485b6ae89f" xmpMM:OriginalDocumentID="xmp.did:77af533c-54fa-f44b-a5a4-7080cd7c6400"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:77af533c-54fa-f44b-a5a4-7080cd7c6400" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:7af6382a-5db8-f840-b3e3-149686d7e425" stEvt:when="2022-09-01T11:00:50+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>$4  �IDATxڵ��O�P �o���nC�L�qQp�?�1f^B$����.��7��ȓ�Չ�Fa��!1����� c[;v9�=��v�݃i��=;���;_��l�(����r�H⧥����kg컵@G�!��yPׁ���S�G"���K���w��'�#�V?#Bv��1�D*�q�0�h�_�\�t:�0R�d���:c�ۛ`�����d2�����)���j���(S��=���,_/�@0��K��u>��45 ��{��
�s�����<Fe-��h���+�n�^������7�>u���!23� �6_(���	MÔ׹��6�W�b���OWo9��H���;>�d�'��sgNQ�隖3��}Z_5W,!��籘x$�FC@�\6>�5B�(�b/�������e�pn"%��]��#_�m~�J��1�-�%����K �k��������{������=�!-
NC(^�q�\*�a[��^j=��cGOt�3��*�2h��D�M��������k��>��iR�J� �5(�Ϟ<��p�t�/���n�j� �F�6���?�b`����)���?h���m�p��p�e<^ۈ���rb��Q���[���+��	�    IEND�B`�  LeftHTop   TPngImageList	Images192Height Width 	PngImages
BackgroundclWindowName&Copy log entries-console window outputPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:45+01:00" xmp:MetadataDate="2022-09-01T11:00:45+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:24444308-3baf-bb40-aac1-f200719333c9" xmpMM:DocumentID="adobe:docid:photoshop:01e673c1-5be5-5040-9100-b3d323c8450c" xmpMM:OriginalDocumentID="xmp.did:91e04cf8-0434-a342-8c33-34c96bbc864f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:91e04cf8-0434-a342-8c33-34c96bbc864f" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:24444308-3baf-bb40-aac1-f200719333c9" stEvt:when="2022-09-01T11:00:45+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>0�J   �IDATx�c���?�@FdL�5���*v�NO>B���vb8 %1�(C��_��������?��:�j���`ؾsɎ��@j_�zM�#��  �D9 d. R�C�OVz2+]B W� �H��"Tw��
< kaEQ �~bB[aE�\@��Vtl�]C [a�����B���*3-	^X�4py � xV�Y�r4�b@� �7TFF��ô�s)�������0�m;�t�@  �����?/    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:48+01:00" xmp:MetadataDate="2022-09-01T11:00:48+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:511b869f-52f9-344f-ba4c-a637b1ad66f2" xmpMM:DocumentID="adobe:docid:photoshop:deddd1a5-dfda-7742-97c1-5094c07dbbf0" xmpMM:OriginalDocumentID="xmp.did:bc5e0618-0e49-9245-9876-d10c035fda57"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:bc5e0618-0e49-9245-9876-d10c035fda57" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:511b869f-52f9-344f-ba4c-a637b1ad66f2" stEvt:when="2022-09-01T11:00:48+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  �IDATx���KSqǿg�M77���Y�i�]0�%],1F��uyt!��2{���B��B�2�nЋ��$��f�ZZkk�1w��r���;�	�|�/�3��������y6��8,��@:��k7���#��y�bV͉G���z��w�`�b2�C
��<�)e0T��W�C���s�݋dx����5��ӗ(p�i�yz W�=��ejA��Y�~��"�o���!i��҆p<!ieyhӪ�X"��`O>�I\
JB^���2	�9�=r��S0�ɥ��u%Ti)~=�ǡ�� ��P���y�p�l_k
�h�ΊY���p,!d����Z%����ṓŹ�ND@��;�`���&Of�!p�iE��@�*l��G����ꆍ p	N0�˜����Q �WO���)�d���K8�|���0���FbB[��?y��!27T�I�k�/U$[�W�}��tLuK_%���6�xC���jz6�f�p{a2R�Q���������*��T��?�$��m�4�"M�YS��M�998��q�h5��_a"m��v^jK��da�̀�]���2��������:X�x5�Gۉ�x)�h�pF��iѵ�<s ^gM�}v�i�0���]C���V�����7�����8�
�h)/����P�4ӤP{����n��J*�@K9���>�yC9��"5������    IEND�B`� 
BackgroundclWindowName"Auto adjust size of console windowPngImage.Data
	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:51+01:00" xmp:MetadataDate="2022-09-01T11:00:51+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:da02287d-009e-b047-8f28-d1aacd00520d" xmpMM:DocumentID="adobe:docid:photoshop:3fee81ce-9a82-8e4d-acb7-0f328a999057" xmpMM:OriginalDocumentID="xmp.did:6740a737-68d9-4f4a-96f7-d113312510c4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:6740a737-68d9-4f4a-96f7-d113312510c4" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:da02287d-009e-b047-8f28-d1aacd00520d" stEvt:when="2022-09-01T11:00:51+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�:�  �IDATx��YkQ�O^��`���҅����nZmҦ|��E�D)m�����Mm�WA)��'�TM7[�""-MR�6��fq�I���L�0/��0�;������sf�l�<� ���u](>7�`��O] �:�D��OWu�~�F�|�M��S��T�d��E�39�qt�����k?V��kH��Û� E
g�8`�Ӂ�_�z]:01w+�(8��ZX�e����}4�܅K��PHZdK����F�e4g��o8{�"�	j"��b Z�o\��V'�3�C#�ԉ�Fp [E�����͠�G�)U��FI�J�B ��~���9?�&���1�j/ �t_���Tk~����Դ���8���@<�Xl��g�P�M�`ǝ�5�0�Vh<���ʧeC��
�@ �%x�j�Vg�ϯ��d�j���gaia��?�Wɝ�1����=�Ym<�z5 �56#ݗ�4<��A2I �[���	4���^Ie,����T%��� ��>X$���d� �X�{��3>�Z˹���kT���Q��;��8 �ZTk^n<�����{G`g0�����`��#���|o�����T� (g�ҁA��˴�݅%���p�� ��B:�" ̬j�K�LF�N>��Pp�M��u�XN�:�t(33T���²��N"�ή��4�O&�! ��T���^��D�]�MOS���L �}j�j/��@�����������W    IEND�B`�  Left�Top     TPF0TCopyDialog
CopyDialogLeftkTop� HelpType	htKeywordHelpKeywordui_copyBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
CopyDialogClientHeight� ClientWidth7Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize7�  
TextHeight TImageImageLeftTopWidth Height AutoSize	  TLabelDirectoryLabelLeft.TopWidth� HeightCaption)Copy 2 selected files to remote directory  THistoryComboBoxLocalDirectoryEditLeft.TopWidth�HeightAutoCompleteAnchorsakLeftakTopakRight DropDownCountTabOrder TextLocalDirectoryEditOnChangeControlChangeOnExitLocalDirectoryEditExit  THistoryComboBoxRemoteDirectoryEditLeft.TopWidthHeightAutoCompleteAnchorsakLeftakTopakRight DropDownCount	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  TButtonOkButtonLeft3Top� WidthPHeightAnchorsakTopakRight CaptionOKDefault	ModalResultTabOrderOnDropDownClickOkButtonDropDownClick  TButtonCancelButtonLeft�Top� WidthPHeightAnchorsakTopakRight Cancel	CaptionAvbrytModalResultTabOrder  TButtonLocalDirectoryBrowseButtonLeft�TopWidthPHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClickLocalDirectoryBrowseButtonClick  	TCheckBoxQueueCheck2Left
TopxWidth=HeightCaption1Transfer in &background (add to transfer queue) XTabOrderOnClickControlChange  TButton
HelpButtonLeft�Top� WidthPHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  	TCheckBoxNeverShowAgainCheckLeft
Top� Width� HeightCaption$   &Visa inte den här dialogrutan igenTabOrder
OnClickNeverShowAgainCheckClick  TButtonTransferSettingsButtonLeftTop� Width� HeightCaption   Överförin&gsinställningar...StylebsSplitButtonTabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxCopyParamGroupLeftTop7Width'Height;AnchorsakLeftakTopakRight Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize';  TLabelCopyParamLabelLeft	TopWidthHeight#AnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamGroupClick   TPanelShortCutHintPanelLeft Top� Width7Height&AlignalBottom
BevelOuterbvNoneParentBackgroundTabOrder	
DesignSize7&  TLabelShortCutHintLabelLeftTopWidth'Height AnchorsakLeftakTopakRightakBottom AutoSizeCaption�   I Commander-gränssnittet används kortkommandot F5 för att överföra filer. Om du vill använda kommandot för att uppdatera en filpanel, klicka här för att gå till inställningar.ShowAccelCharWordWrap	OnClickShortCutHintLabelClick   
TPopupMenuOkMenuLeft�TopE 	TMenuItemDownloadItemCaption
&Ladda nerDefault	OnClickDownloadItemClick  	TMenuItem
BrowseItemCaption	   &BläddraOnClickBrowseItemClick       TPF0TCopyLocalDialogCopyLocalDialogLeft Top HelpType	htKeywordHelpKeywordui_copy_localBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCopyLocalDialogClientHeight~ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�~ 
TextHeight TImageImageLeftTopWidth Height AutoSize	  TLabelDirectoryLabelLeft.TopWidth?HeightCaption   &Målsökväg:FocusControlDirectoryEdit  THistoryComboBoxDirectoryEditLeft.TopWidthsHeightAutoCompleteAnchorsakLeftakTopakRight DropDownCountTabOrder TextDirectoryEditOnExitDirectoryEditExit  TButtonOkButtonLeft� Top7WidthPHeightAnchorsakTopakRight CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftQTop7WidthPHeightAnchorsakTopakRight Cancel	CaptionAvbrytModalResultTabOrder  TButtonLocalDirectoryBrowseButtonLeft�TopWidthPHeightCaption   &Bläddra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButton
HelpButtonLeft�Top7WidthPHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  	TCheckBoxNeverShowAgainCheckLeft
Top;Width� HeightCaption$   &Visa inte den här dialogrutan igenTabOrder  TPanelShortCutHintPanelLeft TopXWidth�Height&AlignalBottom
BevelOuterbvNoneParentBackgroundTabOrder
DesignSize�&  TLabelShortCutHintLabelLeftTopWidth�Height AnchorsakLeftakTopakRightakBottom AutoSizeCaption�   I Commander-gränssnittet används kortkommandot F5 för att överföra filer. Om du vill använda kommandot för att uppdatera en filpanel, klicka här för att gå till inställningar.ShowAccelCharWordWrap	OnClickShortCutHintLabelClick      TPF0TCopyParamCustomDialogCopyParamCustomDialogLeftvTop� HelpType	htKeywordHelpKeywordui_transfer_customBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption   ÖverföringsinställningarClientHeight�ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQuery
DesignSize�� 
TextHeight TButtonOkButtonLeft� Top�WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft$Top�WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  �TCopyParamsFrameCopyParamsFrameLeftTopWidth�Height�HelpType	htKeywordTabOrder   TButton
HelpButtonLeftzTop�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick      TPF0TCopyParamPresetDialogCopyParamPresetDialogLeftTopzHelpType	htKeywordHelpKeywordui_transfer_presetBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCopyParamPresetDialogClientHeight,ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�, 
TextHeight TLabelLabel1LeftTopWidthaHeightCaption   Förinställnings&beskrivningFocusControlDescriptionEdit  TButtonOkButtonLeft�TopWidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft:TopWidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TEditDescriptionEditLeftTopWidth�Height	MaxLength� TabOrder OnChangeControlChange  �TCopyParamsFrameCopyParamsFrameLeftTop2Width�Height�HelpType	htKeywordTabOrder  	TGroupBox	RuleGroupLeft�TopYWidthHeight�AnchorsakLeftakTopakRightakBottom Caption   Regler för automatiskt valTabOrder
DesignSize�  TLabelLabel2Left	TopWidthYHeightCaption   Mask värdna&mnFocusControlHostNameEdit  TLabelLabel3Left	TopEWidthWHeightCaption   Mask an&vändarnamnFocusControlUserNameEdit  TLabelLabel4Left	ToptWidth}HeightCaption   Mask &fjärrkatalogFocusControlRemoteDirectoryEdit  TLabelLabel5Left
Top� WidthpHeightCaptionMask &lokal katalogFocusControlLocalDirectoryEdit  TEditHostNameEditLeft	Top(Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnExitMaskEditExit  TEditUserNameEditLeft	TopWWidth� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditRemoteDirectoryEditLeft	Top� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TEditLocalDirectoryEditLeft	Top� Width� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChangeOnExitMaskEditExit  TButtonCurrentRuleButtonLeft	Top� WidthPHeightCaptionAktuellTabOrderOnClickCurrentRuleButtonClick  TStaticTextRuleMaskHintTextLeft~Top� Width� Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionMasktipsTabOrderTabStop	   	TCheckBoxHasRuleCheckLeft�TopBWidthHeightAnchorsakLeftakTopakRight Caption'   Välj automatiskt förinställning närTabOrderOnClickControlChange  TButton
HelpButtonLeft�TopWidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick     TPF0TCopyParamsFrameCopyParamsFrameLeft Top Width�Height�HelpType	htKeywordFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 
ParentFontTabOrder  	TGroupBoxCommonPropertiesGroupLeft� Top� Width� Height|Caption
AlternativTabOrder
DesignSize� |  TLabelSpeedLabel3Left	Top^WidthFHeightCaption&Hastighet (kB/s)FocusControl
SpeedCombo  	TCheckBoxPreserveTimeCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Behåll tidsstä&mpelParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxCommonCalculateSizeCheckLeftTopDWidth� HeightAnchorsakLeftakTopakRight Caption   B&eräkna total storlekParentShowHintShowHint	TabOrderOnClickControlChange  THistoryComboBox
SpeedComboLeftoTop[WidtheHeightAutoCompleteTabOrderText
SpeedComboOnExitSpeedComboExitItems.Strings	Unlimited10245122561286432168   	TCheckBoxPreserveTimeDirsCheckLeftTop-Width� HeightAnchorsakLeftakTopakRight CaptionInklusive katalogerParentShowHintShowHint	TabOrderOnClickControlChange   	TGroupBoxLocalPropertiesGroupLeft� TopWidth� Height1CaptionNedladdningsalternativTabOrder
DesignSize� 1  	TCheckBoxPreserveReadOnlyCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Behåll skrivsky&ddParentShowHintShowHint	TabOrder    	TGroupBoxRemotePropertiesGroupLeftTop� Width� Height� Caption   ÖverföringsalternativTabOrder 	TCheckBoxPreserveRightsCheckLeftTopWidth� HeightCaption   Sätt fil&rättigheterParentShowHintShowHint	TabOrder OnClickControlChange  
TComboEdit
RightsEditLeftTop-Width{Height
ButtonHint   Konfigurera filrättigheterClickKey@ParentShowHintShowHint	TabOrderText
RightsEditOnButtonClickRightsEditButtonClickOnExitRightsEditExitOnContextPopupRightsEditContextPopup  	TCheckBoxIgnorePermErrorsCheckLeftTopHWidth� HeightCaption   Ign&orera filrättighetsfelParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxClearArchiveCheckLeftTop_Width� HeightCaptionRensa 'Arki&v' attributTabOrder  	TCheckBoxRemoveCtrlZAndBOMCheckLeftTopvWidth� HeightCaptionRemo&ve BOM and EOF marks XTabOrderOnClickControlChange  	TCheckBoxEncryptNewFilesCheckLeftTop� Width� HeightCaption&Kryptera nya filerTabOrderOnClickControlChange   	TGroupBoxChangeCaseGroupLeft"TopWidth� Height� Caption   Ändra filnamnTabOrder
DesignSize� �   TRadioButtonCCLowerCaseShortButtonLeftTop[Width� HeightAnchorsakLeftakTopakRight CaptionGemener &8.3TabOrder  TRadioButtonCCNoChangeButtonLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   I&ngen förändringTabOrder   TRadioButtonCCUpperCaseButtonLeftTop-Width� HeightAnchorsakLeftakTopakRight Caption	&VersalerTabOrder  TRadioButtonCCLowerCaseButtonLeftTopDWidth� HeightAnchorsakLeftakTopakRight Caption&GemenerTabOrder  	TCheckBoxReplaceInvalidCharsCheckLeftToprWidth� HeightCaption   &Ersätt '\:*?' ...TabOrderOnClickControlChange   	TGroupBoxTransferModeGroupLeftTopWidthHeight� Caption   ÖverföringslägeTabOrder 
DesignSize�   TLabelAsciiFileMaskLabelLeft	Top[Width� HeightAnchorsakLeftakTopakRight Caption'   Överför följande &filer i textläge:FocusControlAsciiFileMaskCombo  TRadioButtonTMTextButtonLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption&Text (text, html, skript, ...)TabOrder OnClickControlChange  TRadioButtonTMBinaryButtonLeftTop-Width� HeightAnchorsakLeftakTopakRight Caption   &Binärt (arkiv, doc, ...)TabOrderOnClickControlChange  TRadioButtonTMAutomaticButtonLeftTopDWidth� HeightAnchorsakLeftakTopakRight Caption&AutomatisktTabOrderOnClickControlChange  THistoryComboBoxAsciiFileMaskComboLeft	TopmWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextAsciiFileMaskComboOnExitValidateMaskComboExit   	TGroupBox
OtherGroupLeftTopPWidth�Height� Caption   ÖvrigtTabOrder
DesignSize��   TLabelIncludeFileMaskLabelLeft	TopWidth4HeightCaptionFilmas&kFocusControlIncludeFileMaskCombo  THistoryComboBoxIncludeFileMaskComboLeft	Top(WidthZHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextIncludeFileMaskComboOnExitValidateMaskComboExit  TButtonIncludeFileMaskButtonLeftiTop'WidthPHeightAnchorsakTopakRight Caption&Redigera...TabOrderOnClickIncludeFileMaskButtonClick  	TCheckBoxNewerOnlyCheckLeftTopQWidth� HeightCaption!Endast &nya och uppdaterade filerParentShowHintShowHint	TabOrderOnClickControlChange  TStaticTextIncludeFileMaskHintTextLeft� Top?Width}Height	AlignmenttaRightJustifyAutoSizeCaptionmasktipsTabOrderTabStop	  	TCheckBoxExcludeHiddenFilesCheckLeft� TopQWidth� HeightCaptionExkludera &dolda filerParentShowHintShowHint	TabOrderOnClickControlChange  	TCheckBoxExcludeEmptyDirectoriesCheckLeftTophWidth� HeightCaptionE&xkludera tomma katalogerParentShowHintShowHint	TabOrderOnClickControlChange       TPF0TCreateDirectoryDialogCreateDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeywordui_create_directoryBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSkapa katalogClientHeightClientWidthQColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizeQ 
TextHeight TLabel	EditLabelLeftTopWidth^HeightCaptionNytt &katalognamn:FocusControlDirectoryEdit  TEditDirectoryEditLeftTopWidthAHeightAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextDirectoryEditOnChangeDirectoryEditChange  TPanel	MorePanelLeft Top2WidthQHeight� AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder
DesignSizeQ�   	TGroupBoxAttributesGroupLeftTopWidthAHeight� AnchorsakLeftakTopakRightakBottom Caption
EgenskaperTabOrder  �TRightsFrameRightsFrameLeftTop'WidthHeightbTabOrder �	TCheckBoxDirectoriesXCheckVisible   	TCheckBoxSetRightsCheckLeftTopWidth� HeightCaption   Sätt fil&rättigheterParentShowHintShowHint	TabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeftTop� Width-HeightCaption*   Använd &samma inställningar nästa gångTabOrder    TButtonOKBtnLeftMTop� WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft� Top� WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft� Top� WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick      TPF0TCustomCommandDialogCustomCommandDialogLeft�Top� HelpType	htKeywordHelpKeywordui_customcommandBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionCustomCommandDialogClientHeightClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize� 
TextHeight 	TGroupBoxGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight TabOrder 
DesignSize��   TLabelDescriptionLabelLeft	Top	Width?HeightCaption&BeskrivningFocusControlDescriptionEdit  TLabelLabel1Left	Top8WidthgHeightCaption&Eget kommando:FocusControlCommandEdit  TLabelShortCutLabelLeft	Top� WidthdHeightCaptionKor&tkommando:FocusControlShortCutCombo  TEditDescriptionEditLeft	TopWidth�HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  THistoryComboBoxCommandEditLeft	TopJWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength TabOrderOnChangeControlChange	OnGetDataCommandEditGetData	OnSetDataCommandEditSetData  	TCheckBoxApplyToDirectoriesCheckLeftTop� Width� HeightCaption   &Tillämpa på katalogerTabOrderOnClickControlChange  	TCheckBoxRecursiveCheckLeft� Top� Width� HeightCaption   Kör &rekursivtTabOrderOnClickControlChange  TRadioButtonLocalCommandButtonLeft� TopsWidth� HeightCaption&Lokalt kommandoTabOrderOnClickControlChange  TRadioButtonRemoteCommandButtonLeftTopsWidth� HeightCaption   &FjärrkommandoTabOrderOnClickControlChange  	TCheckBoxShowResultsCheckLeftTop� Width� HeightCaption!   &Visa resultat i terminalfönsterTabOrderOnClickControlChange  	TCheckBoxCopyResultsCheckLeftTop� Width� HeightCaption&Kopiera resultat till urklippTabOrder	OnClickControlChange  TStaticTextHintTextLeftATopaWidthvHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  	TComboBoxShortCutComboLeft� Top� Width� HeightTabOrder
  	TCheckBoxRemoteFilesCheckLeft� Top� Width� HeightCaption   &Använd fjärrfilerTabOrderOnClickControlChange   TButtonOkButtonLeft� Top� WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft"Top� WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftxTop� WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPF0TCustomDialogCustomDialogLeft�Top� BorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSave session as siteXClientHeight*ClientWidthjColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenter
DesignSizej* 
TextHeight TButtonOKButtonLeftfTop	WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top	WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder   TButton
HelpButtonLeftTop	WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TPF0TCustomScpExplorerFormCustomScpExplorerFormLeft� Top� CaptionCustomScpExplorerFormClientHeight�ClientWidth`Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 
KeyPreview	OnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnClose	FormCloseOnCloseQueryFormCloseQueryOnConstrainedResizeFormConstrainedResizeOnShowFormShow
TextHeight 	TSplitterQueueSplitterLeft TopWidth`HeightCursorcrSizeNSHintR   Dra för att ändra storlek på kölistan. Dubbelklicka för att dölja kölistan.AlignalBottomAutoSnapMinSizeFResizeStylersUpdateOnCanResizeQueueSplitterCanResize  TTBXDockTopDockLeft Top Width`Height	FixAlign	  TPanelRemotePanelLeft Top'Width`Height� AlignalClient
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder  	TSplitterRemotePanelSplitterLeft� Top Height� CursorcrSizeWEAutoSnapMinSizeFResizeStylersUpdate  TTBXStatusBarRemoteStatusBarLeft Top� Width`HeightPanels ParentShowHintShowHint	UseSystemFontOnClickRemoteStatusBarClickOnMouseDownRemoteStatusBarMouseDown  TPanelRemoteDirPanelLeft� Top Width�Height� AlignalClient
BevelOuterbvNoneTabOrder TUnixDirViewRemoteDirViewLeft Top Width�Height� AlignalClientDoubleBuffered	FullDrag	HideSelectionIconOptions.AutoArrange	ParentDoubleBuffered	PopupMenu&NonVisualDataModule.RemoteDirViewPopupTabOrder OnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterRemoteDirViewEnterOnExitDirViewExit	OnKeyDownDirViewKeyDown
OnKeyPressDirViewKeyPressOnResizeRemoteDirViewResize
NortonLikenlOffUnixColProperties.ExtWidthUnixColProperties.TypeVisibleOnDDDragFileNameRemoteFileControlDDDragFileNameOnBusyDirViewBusyOnChangeFocusDirViewChangeFocusOnSelectItemDirViewSelectItemOnStartLoadingRemoteDirViewStartLoadingOnLoadedDirViewLoaded
OnExecFileDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayDirViewGetOverlayOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDDragDetectRemoteFileControlDDDragDetectOnDDEndRemoteFileControlDDEndOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectOnContextPopupRemoteDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnDisplayPropertiesRemoteDirViewDisplayPropertiesDirViewStyle	dvsReportOnReadRemoteDirViewReadOnStartReadingRemoteDirViewStartReadingOnThumbnailNeededRemoteDirViewThumbnailNeeded  TTBXToolbarReconnectToolbarLeft� ToppWidthkHeightCaptionReconnectToolbarImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem254Action*NonVisualDataModule.ReconnectSessionAction    TPanelRemoteDrivePanelLeft Top Width� Height� AlignalLeft
BevelOuterbvNoneTabOrder TUnixDriveViewRemoteDriveViewLeft Top Width� Height� DirViewRemoteDirViewOnDDDragFileNameRemoteFileControlDDDragFileNameOnDDEndRemoteFileControlDDEndUseSystemContextMenuOnDDDragEnterFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDQueryContinueDrag$RemoteFileControlDDQueryContinueDragOnDDChooseEffectRemoteFileContolDDChooseEffectOnDDGiveFeedbackRemoteFileControlDDGiveFeedbackOnDDDragDetectRemoteFileControlDDDragDetectOnDDFileOperation RemoteFileControlDDFileOperationOnDDCreateDragFileList%RemoteFileControlDDCreateDragFileListOnDDCreateDataObject#RemoteFileControlDDCreateDataObjectAlignalClientDoubleBuffered	HideSelectionIndentParentColorParentDoubleBufferedReadOnly	TabOrder OnEnterRemoteDriveViewEnterOnBusyDirViewBusy    TPanel
QueuePanelLeft Top!Width`Height� AlignalBottom
BevelOuterbvNoneTabOrder 
TPathLabel
QueueLabelLeft Top WidthlHeightIndentVerticalAutoSizeVertical	OnGetStatusQueueLabelGetStatusAutoSizeTransparent  	TSplitterQueueFileListSplitterLeft TopuWidthlHeightCursorcrSizeNSHintd   Dra för att ändra storlek på köfilens lista. Dubbelklicka för att dölja listan över köfiler.AlignalBottomAutoSnapMinSize
ResizeStylersUpdateOnCanResizeQueueFileListSplitterCanResize  	TListView
QueueView3Left Top/WidthlHeightFAlignalClientColumnsCaption	OperationMinWidthWidthF Caption   KällaMinWidthWidth�  Caption   MålMinWidthWidth�  	AlignmenttaRightJustifyCaption
   ÖverförtMinWidthWidthP 	AlignmenttaRightJustifyCaptionTidMinWidthWidthP 	AlignmenttaRightJustifyCaption	HastighetMinWidthWidthP 	AlignmenttaCenterCaption
UtvecklingMinWidthWidthP  ColumnClickDoubleBuffered	DragModedmAutomaticReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuNonVisualDataModule.QueuePopupSmallImagesGlyphsModule.QueueImagesStateImagesGlyphsModule.QueueImagesTabOrder 	ViewStylevsReportOnChangeQueueView3ChangeOnContextPopupQueueView3ContextPopup
OnDeletionQueueView3Deletion	OnEndDragQueueView3EndDragOnEnterQueueView3EnterOnExitQueueView3Exit
OnDragDropQueueView3DragDrop
OnDragOverQueueView3DragOverOnSelectItemQueueView3SelectItemOnStartDragQueueView3StartDrag  TTBXDock	QueueDockTagLeft TopWidthlHeight	AllowDrag TTBXToolbarQueueToolbarLeft Top CaptionQueueToolbarImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder  TTBXItemQueueEnableItemAction%NonVisualDataModule.QueueEnableAction  TTBXSeparatorItemTBXSeparatorItem203  TTBXItem
TBXItem201Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem
TBXItem202Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem
TBXItem203Action)NonVisualDataModule.QueueItemPromptAction  TTBXItem
TBXItem204Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem195Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem194Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem
TBXItem205Action)NonVisualDataModule.QueueItemDeleteAction  TTBXSeparatorItemTBXSeparatorItem201  TTBXItem
TBXItem206Action%NonVisualDataModule.QueueItemUpAction  TTBXItem
TBXItem207Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem57  TTBXItem"QueueDeleteAllDoneQueueToolbarItemAction,NonVisualDataModule.QueueDeleteAllDoneAction  TTBXSeparatorItemTBXSeparatorItem202  TTBXSubmenuItemTBXSubmenuItem27Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem211Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem225Action3NonVisualDataModule.QueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem173Action0NonVisualDataModule.QueueSuspendOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem226Action1NonVisualDataModule.QueueShutDownOnceEmptyAction2	RadioItem	   TTBXItem
TBXItem208Action*NonVisualDataModule.QueuePreferencesAction    	TListViewQueueFileListLeft TopxWidthlHeightAlignalBottomColumns  DoubleBuffered		OwnerData	ReadOnly	ParentDoubleBufferedShowColumnHeadersTabOrderTabStop	ViewStylevsReportOnCustomDrawItemQueueFileListCustomDrawItemOnDataQueueFileListDataOnEnterQueueFileListEnterExitOnExitQueueFileListEnterExitOnResizeQueueFileListResize   TThemePageControlSessionsPageControlLeft TopWidth`Height
ActivePage	TabSheet1AlignalTopDoubleBuffered	ParentDoubleBufferedParentShowHintShowHint	TabOrderTabStopOnChangeSessionsPageControlChangeOnContextPopupSessionsPageControlContextPopup
OnDragDropSessionsPageControlDragDrop
OnDragOverSessionsPageControlDragOverOnMouseDownSessionsPageControlMouseDownOnResizeSessionsPageControlResizeOnTabButtonClick!SessionsPageControlTabButtonClick	OnTabHintSessionsPageControlTabHint TThemeTabSheet	TabSheet1Caption	TabSheet1   TTBXDockMessageDockTagLeft Top	Width`Height		AllowDragFixAlign	VisibleOnRequestDockMessageDockRequestDock  TApplicationEventsApplicationEventsOnDeactivateApplicationEventsDeactivate
OnMinimizeApplicationMinimizeOnModalBeginApplicationEventsModalBegin	OnRestoreApplicationRestoreLeftXTop�     TPF0TEditMaskDialogEditMaskDialogLeftqTopHelpType	htKeywordHelpKeywordui_editmaskBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRedigera filmaskClientHeightClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 
KeyPreview	PositionpoOwnerFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize� 
TextHeight 	TGroupBox
FilesGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption	FilmaskerTabOrder 
DesignSize��   TLabelLabel3Left	TopWidthBHeightCaption&Inkludera filer:FocusControlIncludeFileMasksMemo  TLabelLabel1Left� TopWidthCHeightCaption&Exkludera filer:FocusControlExcludeFileMasksMemo  TMemoIncludeFileMasksMemoLeft	Top(Width� Height� AnchorsakLeftakTopakBottom Lines.StringsIncludeFileMasksMemo 
ScrollBars
ssVerticalTabOrder OnChangeControlChangeOnExitFileMasksMemoExit  TMemoExcludeFileMasksMemoLeft� Top(Width� Height� AnchorsakLeftakTopakBottom Lines.StringsExcludeFileMasksMemo 
ScrollBars
ssVerticalTabOrderOnChangeControlChangeOnExitFileMasksMemoExit   TButtonOKBtnLeft� Top�WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft,Top�WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeft�Top�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClearButtonLeft� Top�WidthPHeightAnchorsakRightakBottom Caption&RensaTabOrderOnClickClearButtonClick  	TGroupBoxDirectoriesGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight CaptionKatalogmaskerTabOrder
DesignSize��   TLabelLabel2Left	TopWidthdHeightCaptionI&nkludera kataloger:FocusControlIncludeDirectoryMasksMemo  TLabelLabel4Left� TopWidtheHeightCaptionE&xkludera kataloger:FocusControlExcludeDirectoryMasksMemo  TMemoIncludeDirectoryMasksMemoLeft	Top(Width� HeightsAnchorsakLeftakTopakBottom Lines.StringsIncludeDirectoryMasksMemo 
ScrollBars
ssVerticalTabOrder OnChangeControlChangeOnExitDirectoryMasksMemoExit  TMemoExcludeDirectoryMasksMemoLeft� Top(Width� HeightsAnchorsakLeftakTopakBottom Lines.StringsExcludeDirectoryMasksMemo 
ScrollBars
ssVerticalTabOrderOnChangeExcludeDirectoryMasksMemoChangeOnExitDirectoryMasksMemoExit  	TCheckBoxExcludeDirectoryAllCheckLeft� Top� Width� HeightAnchorsakLeftakBottom Caption&Alla (rekursera inte)TabOrderOnClickExcludeDirectoryAllCheckClick   	TGroupBox	MaskGroupLeftTop�Width�HeightYAnchorsakLeftakTopakRight CaptionMaskTabOrder
DesignSize�Y  TMemoMaskMemoLeft	TopWidth�Height:TabStopAnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneLines.StringsMaskMemo 
ScrollBars
ssVerticalTabOrder    TStaticTextMaskHintTextLeftQTop�Width� Height	AlignmenttaRightJustifyAutoSizeCaptionmasktipsTabOrderTabStop	    TPF0TEditorForm
EditorFormLeft;Top� HelpType	htKeywordHelpKeyword	ui_editorBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp Caption
EditorFormClientHeight}ClientWidthaColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 	Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ��������������������������������������������������������������������Leo�t�����������������������������������������������������������������������������������������������������������                                                                            ��������������������������������������������������������������������k���OKG�Kak�����������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������OKG�OKG�LML�t�����������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������KOO�OKG�OKG�OKG�Gv������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������Ojv�OKG�NLI�&i�� ���	���������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������}���ERW�y�� ��� ��� ��� ���C�������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������� ��� ��� ��� ��� ��� ������������������������������������������������������������������������������                                                                            ����������������������������������������������������������������������������!��� ��� ��� ��� ��� ��� ��� ��� ���J�������������������������������������������������������������������                                                                            ����������������������������������������������������������������������������f��� ��� ��� ��� ��� ��� ��� ��� ������s���������������������������������������������������������������                                                                            �������������������������������������������������������������������������������� ��� ��� ��� ��� ��� ��� ���	���������������������������������������������������������������������                                                                            ����������������������������������������������������������������������������������� ��� ��� ��� ������������������)�����������������������������������������������������������                                                                            ��������������������������������������������������������������������������������3��� ��� ������#���%���#��� ������������V�������������������������������������������������������                                                                            ��������������������������������������������������������������������������������w��� ��� ������+���(���%���#��� ����������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������*������-���.���+���(���%���"���������������������������������������������������������������                                                                            ����������������������������������������������������������������������������������������5���2���0���-���*���'���$���!������������9�����������������������������������������������                                                                            ��������������������������������������������������������������������������������������������5���2���/���,���)���&���#��� ������������o�������������������������������������������                                                                            ��������������������������������������������������������������������������������������������T���4���1���.���+���(���%���"�������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������:���3���0���-���*���'���$���!������������(���������������������������������������                                                                            ����������������������������������������������������������������������������������������������������5���2���/���,���)���&���#���!������������N�����������������������������������                                                                            ����������������������������������������������������������������������������������������������������l���4���1���.���,���(���&���#��� ��������������������������������������������                                                                            ��������������������������������������������������������������������������������������������������������E���3���0���.���+���(���%���"�������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������5���3���0���-���*���'���$���!������������6���������������������������                                                                            ����������������������������������������������������������������������������������������������������������������5���2���/���,���)���&���#��� ������������l�����������������������                                                                            ����������������������������������������������������������������������������������������������������������������U���4���1���.���+���(���%���"�����������������������������������                                                                            ��������������������������������������������������������������������������������������������������������������������<���3���0���-���*���'���$���"������������&�������������������                                                                            ������������������������������������������������������������������������������������������������������������������������5���2���/���,���)���&���$���!������������J���������������                                                                            ������������������������������������������������������������������������������������������������������������������������n���4���1���/���,���(���&���#��� ������������������������                                                                            ����������������������������������������������������������������������������������������������������������������������������H���3���1���.���+���(���%���"�����������������������                                                                            ��������������������������������������������������������������������������������������������������������������������������������7���3���0���-���*���'���$���!������������2�������                                                                            ������������������������������������������������������������������������������������������������������������������������������������5���2���/���,���)���&���#��� ������������F���                                                                            ������������������������������������������������������������������������������������������������������������������������������������X���4���1���.���+���(���%���"�����������������_                                                                        ����������������������������������������������������������������������������������������������������������������������������������������=���3���0���-���*���'���$���"�����������������$                                                                    ��������������������������������������������������������������������������������������������������������������������������������������������5���2���/���,���)���'���$���!��������������� ��                                                                ��������������������������������������������������������������������������������������������������������������������������������������������V���4���2���/���,���)���&���#��� ���������������                                                                ������������������������������������������������������������������������������������������������������������������������������������������������H���4���1���.���+���(���%���"������������h��·��@                                                            ����������������������������������������������������������������������������������������������������������������������������������������������������7���3���0���-���*���'���$���!���(����ǻ������寯�                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������5���2���/���,���)���&���W��������ÿ�������������                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������_���4���1���.���.����������������������������������m                                                    ������������������������������������������������������������������������������������������������������������������������������������������������������������:���3���L���������������������������¿������f~�� 9�$                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������T�ޅ������������������������������������9b��=��<�� +�                                            �����������������������������������������������������������������������������������������������������������������������������������������������������������<    ��������������������������������M��=��=��=��=؋                                            �������������������������������������������������������������������������������������������������������������������������������������������������������<        �����������������������n���P��G��?��=��=��<�� <�H                                        ���������������������������������������������������������������������������������������������������������������������������������������������������<                ���;������������E|��\��T��M��	E��=��=��=��=�� 3�                                    �����������������������������������������������������������������������������������������������������������������������������������������������<                        ��������*k��$g�� b��Z��R��K��C��=��=��=��<٩                                    �������������������������������������������������������������������������������������������������������������������������������������������<                              �#f��$g��$g��$g��`��X��P��H��@��=��=��=��                                    ���������������������������������������������������������������������������������������������������������������������������������������<                                    #c�$$g��$g��$g��"e��]��V��N��
F��>��=��=ج                                    �����������������������������������������������������������������������������������������������������������������������������������<                                            $e�]$g��$g��$g��!c��[��S��L��D��<ٚ 3�
                                    �������������������������������������������������������������������������������������������������������������������������������<                                                    $g�$g��$g��$g��a��Y��Q��H�Q                                                                                                                                                                                                                                [�#g��$g��$g��#f��^�N�                                                                                                                                                                                                                                        "f�-#f��$g��#f�v  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ���������������������������������     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��      ��      ��      �      ?�      �     �     �     �    ? �     �    ���   ���   ���������?�������������������������������(   0   `          �%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ������������������������������������������������������������������������������������������������������������������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            ��������������������������������������������������������z���������������������������������������������������������������������������                                                            ��������������������������������������������������������LML�Lcm���������������������������������������������������������������������                                                            ��������������������������������������������������������Kcm�OKG�KNN�|���������������������������������������������������������������                                                            ��������������������������������������������������������o���OKG�NKH�(h��C�����������������������������������������������������������                                                            ������������������������������������������������������������ERV�x�� ��� ����������������������������������������������������������                                                            ��������������������������������������������������������������� ��� ��� ��� ��� ���C�����������������������������������������������                                                            ������������������������������������������������������������X��� ��� ��� ��� ��� ��� ���)�������������������������������������������                                                            ���������������������������������������������������������������� ��� ��� ��� ��� ���������L���������������������������������������                                                            ���������������������������������������������������������������� ��� ��� ������������������������������������������������������                                                            ����������������������������������������������������������������-��� ������*���&���"��������������������������������������������                                                            ����������������������������������������������������������������{���������,���)���%���!���������4�������������������������������                                                            ��������������������������������������������������������������������_���3���/���+���(���$��� ���������j���������������������������                                                            ������������������������������������������������������������������������A���2���.���*���&���#������������������������������������                                                            ����������������������������������������������������������������������������5���1���-���)���%���"���������&�����������������������                                                            ����������������������������������������������������������������������������}���4���0���,���(���$���!���������H�������������������                                                            ��������������������������������������������������������������������������������M���2���/���+���'���#����������������������������                                                            ������������������������������������������������������������������������������������6���1���.���*���&���"������������������������                                                            ����������������������������������������������������������������������������������������4���0���,���)���%���!���������1�����������                                                            ����������������������������������������������������������������������������������������b���3���/���,���(���$��� ���������a�������                                                            ��������������������������������������������������������������������������������������������A���2���.���*���'���#������������k���                                                            ������������������������������������������������������������������������������������������������5���1���-���)���%���"��������������$                                                        ����������������������������������������������������������������������������������������������������4���0���,���(���$���!������������ ��                                                    ����������������������������������������������������������������������������������������������������Q���2���/���+���'���#��� ������������                                                    ��������������������������������������������������������������������������������������������������������8���2���.���*���&���"��������������F                                                ������������������������������������������������������������������������������������������������������������4���0���-���)���%���!��������������                                            ������������������������������������������������������������������������������������������������������������h���3���/���,���(���$��� ������������                                            ����������������������������������������������������������������������������������������������������������������<���2���.���*���'���#������������(��e                                        ��������������������������������������������������������������������������������������������������������������������5���1���-���)���%���"������p��¸��쳳�(                                    ��������������������������������������������������������������������������������������������������������������������{���4���0���,���(���0�������¾��������Ӫ��                                ������������������������������������������������������������������������������������������������������������������������:���3���/���g���������������ÿ����������                                �����������������������������������������������������������������������������������������������������������������������<5��07�������������������������������%S�� <�H                            �������������������������������������������������������������������������������������������������������������������<        ���l������������������������
B��=��=�� 5�                        ���������������������������������������������������������������������������������������������������������������<            �������������������V���L��B��=��=��<ٷ                        �����������������������������������������������������������������������������������������������������������<                    �����������8t��^��T��J��?��=��=��<�o                    �������������������������������������������������������������������������������������������������������<                            }��\%h��$g��"e��[��Q��G��=��=��<��                    ���������������������������������������������������������������������������������������������������<                                    $f�$g��$g�� b��X��N��D��=��<ٻ                                                                                                                                                             `�$g��$g��$g��_��U��K��A۞ 3�
                                                                                                                                                                #c�,$g��$g��#f��\��P�S                                                                                                                                                                            $e�]$g��$g�a�                                                                                                                                                                                                                    ������  ������  ������  ������  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �    �  �    �  �      �    ?  �      �      �      �   �  �  �  �  �  �  �  �  �  �����  �����  �����  ������  (   (   P          @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ������������������������������������������������������������������������������������������������������������                                                    ������������������������������������������������������������������������������������������������������������                                                    ��������������������������������������������j���������������������������������������������������������������                                                    ��������������������������������������������o���LML�t�������������������������������������������������������                                                    ������������������������������������������������OKG�OKG�Im~�������������������������������������������������                                                    ������������������������������������������������JPQ�1`w����	�����������������������������������������������                                                    ������������������������������������������������U��� ��� ��� ��� ���C���������������������������������������                                                    ���������������������������������������������������� ��� ��� ��� ��� ���'�����������������������������������                                                    ���������������������������������������������������� ��� ��� ��� ��� ������@�������������������������������                                                    ����������������������������������������������������%��� ������������������~���������������������������                                                    ����������������������������������������������������d��� ��� ���)���%���!���������������������������������                                                    ��������������������������������������������������������A���0���-���(���$���������/�����������������������                                                    ������������������������������������������������������������4���0���,���'���"���������Y�������������������                                                    ����������������������������������������������������������������3���/���*���&���!�������������������������                                                    ����������������������������������������������������������������X���2���-���)���$��� ���������������������                                                    ��������������������������������������������������������������������;���1���,���(���#���������=�����������                                                    ������������������������������������������������������������������������4���/���+���&���"���������v�������                                                    ������������������������������������������������������������������������r���2���.���*���%���!���������u���                                                    ����������������������������������������������������������������������������H���1���-���(���$���������#�����                                                ��������������������������������������������������������������������������������6���0���,���'���"������������ ��                                            ������������������������������������������������������������������������������������3���/���*���&���!�����������t                                            ������������������������������������������������������������������������������������_���2���-���)���%��� �����������5                                        ����������������������������������������������������������������������������������������<���1���,���(���#��������������
                                    ��������������������������������������������������������������������������������������������4���/���+���&���"������������                                    ��������������������������������������������������������������������������������������������x���3���.���*���%���!���������U��K                                ������������������������������������������������������������������������������������������������K���1���-���(���$���(����Ź��ﱱ�                            ����������������������������������������������������������������������������������������������������6���0���,���U����������������������                        ����������������������������������������������������������������������������������������������������h���4��������������������¾�����+W�~                        �������������������������������������������������������������������������������������������������������?������������������������D��=�� :�5                    ���������������������������������������������������������������������������������������������������<    ���"������������^���K��?��=��=�� 7�                �����������������������������������������������������������������������������������������������<            ���b����>x��_��S��G��=��=��<؞                �������������������������������������������������������������������������������������������<                    'j�$g��$g��[��P��D��=��<��                ���������������������������������������������������������������������������������������<                        [�#g��$g��"d��X��L��@��=�`                �����������������������������������������������������������������������������������<                                $g�9$g��$g��a��U��H�.                                                                                                                                            #f�n$g��#f� @�                                                                                                                                                                            �����   �����   �����   �����   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �   �   �   �   �      �   ?   �   ?   �      �      �      �      �      �     �     �  >   �  ~   �  �   �����   �����   (       @          �                                                                                                                                                                                                                                                                                                  ��������������������������������������������������������������������������������������������                                    ��������������������������������������������������������������������������������������������                                    ��������������������������������������������������������������������������������������������                                    ������������������������������������OKG�Ojv�������������������������������������������������                                    ������������������������������������IY`�:Zi������������������������������������������������                                    ������������������������������������k��� ��� ��� ���Q���������������������������������������                                    ���������������������������������������� ��� ��� ��� ���7�����������������������������������                                    ������������������������������������������� ���
���������m�������������������������������                                    ����������������������������������������7������*���$�������������������������������������                                    ��������������������������������������������1���.���(���#������&���������������������������                                    ������������������������������������������������2���,���'���!������L�����������������������                                    ������������������������������������������������b���1���+���%�����������������������������                                    ����������������������������������������������������@���/���)���$�������������������������                                    ��������������������������������������������������������3���-���(���"������4���������������                                    ������������������������������������������������������������2���,���&��� ������j�����������                                    ������������������������������������������������������������Q���0���*���$�����������������                                    ����������������������������������������������������������������8���.���(���#������&�������                                    ��������������������������������������������������������������������2���-���'���!������5��� ��                                ��������������������������������������������������������������������i���1���+���%������������                                ������������������������������������������������������������������������A���/���)���$���������;��8                            ������������������������������������������������������������������������~���3���-���(���)����������⯯�                        ��������������������������������������������������������������������������������2���Y�������������������                        ����������������������������������������������������������������������������������������������������#R��<�a                    �����������������������������������������������������������������������������������a������������N��=��<�� 9�$                �������������������������������������������������������������������������������<    ����c���!c��T��	E��=��=��                ���������������������������������������������������������������������������<          �#g�$g��_��P��A��<��                �����������������������������������������������������������������������<                 `�$g��$g��[��L� 7�                �������������������������������������������������������������������<                        "e�D$g��"d�a                                                                                                                                                                                                                                                                        ���������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �   �  �� �� �� ���������(      0          `	                                                                                                                                                                                                                              ��������������������������������������������������������������������                            ��������������������������������������������������������������������                            ������������������������^}������������������������������������������                            ������������������������Ojv�GV[�������������������������������������                            ����������������������������}�� ���a�������������������������������                            ���������������������������� ��� ��� ���:���������������������������                            ����������������������������!������������o�����������������������                            ����������������������������y���%���)���"��������������������������                            ��������������������������������_���.���'������(�������������������                            ������������������������������������?���,���%������N���������������                            ����������������������������������������2���*���#������������������                            ����������������������������������������}���/���(���!��������������                            ��������������������������������������������L���-���&������8�������                            ������������������������������������������������6���+���$������J���                            ������������������������������������������������k���1���)���"��������[                        ����������������������������������������������������b���/���'��� ������j��                    ��������������������������������������������������������9���,���6�����̸��ƀ��                ��������������������������������������������������������X�݀y���������������0[̈́                �������������������������������������������������������<    ������������N��<�� :�9            ���������������������������������������������������<        �������#e��R��>��=��                                                                            "e�5$g��`��L��<ډ                                                                                #f�n$g��Y�M    ��� ��� �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � @ � � ��� ��� (      (          �                                                                                                          ������������������������������������������������������������                    ������������������������������������������������������������                    ������������������������������������������������������������                    ������������������������^|����������������������������������                    ������������������������Qo}�-u������������������������������                    ���������������������������� ��� ���h�����������������������                    ���������������������������� ���#��������������������������                    ����������������������������P���,���#���!�������������������                    ��������������������������������A���*���!���@���������������                    ������������������������������������0���'������{�����������                    ����������������������������������������.���%��������������                    ����������������������������������������S���+���"���/�������                    ��������������������������������������������6���(������?���                    ��������������������������������������������p���/���&��������r                ������������������������������������������������g���-���>��괻�ϴ��,            ����������������������������������������������������������������Oo��  �        �����������������������������������������������󝙕<���H����8l��=��<ؘ        �����������������������������������������������<        )j�$g��N��=��                                                                 `�$g��_� 7���� � p � p � p � p � p � p � p � p � p � p � p � p � p � 0 �  �   �   �  ��  (                 @                                                                                          ������������������������������������������������                ������������������������������������������������                ����������������(h��[���������������������������                ������������������� ���8�����������������������                ����������������b���'������a�������������������                ��������������������E���(����������������������                ������������������������1���%���#���������������                ����������������������������-���"���D�����������                ����������������������������V���*��������������                ��������������������������������7���'������x���                ��������������������������������u���.���$���9������            ������������������������������������l���q��������            ���������������������������������������������I��=�i        ���������������������������������������<t��Q$g��P��=��                                                    $f�"c��D�)��  �  �  �  �  �  �  �  �  �  �  �  �  �   �   ��  
KeyPreview	OnClose	FormCloseOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
TextHeight TTBXDockTopDockLeft Top WidthaHeight	AllowDrag TTBXToolbarToolBarLeft Top CaptionToolBarImagesEditorImagesOptionstboShowHint ParentShowHintShowHint	TabOrder  TTBXItemTBXItem2Action
SaveAction  TTBXItemTBXItem1ActionSaveAllAction2  TTBXItem	TBXItem16ActionReloadAction  TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem3ActionEditCopy  TTBXItemTBXItem4ActionEditCut  TTBXItemTBXItem5Action	EditPaste  TTBXItemTBXItem6Action
EditDelete  TTBXItemTBXItem7ActionEditSelectAll  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem8ActionEditUndo  TTBXItem	TBXItem17ActionEditRedo  TTBXSeparatorItemTBXSeparatorItem3  TTBXItemTBXItem9Action
FindAction  TTBXItem	TBXItem10ActionReplaceAction  TTBXItem	TBXItem11ActionFindNextAction  TTBXItem	TBXItem12ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemEncodingCaptionKodningHint   Ändra filkodningOptionstboDropdownArrow  TTBXItemDefaultEncodingActionDefaultEncodingAction	RadioItem	  TTBXItemUTF8EncodingActionUTF8EncodingAction	RadioItem	   TTBXColorItem	ColorItemActionColorActionOptionstboDropdownArrow   TTBXItem	TBXItem13ActionPreferencesAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem14Action
HelpAction    TTBXStatusBar	StatusBarLeft TopgWidthaPanelsCaptionLine: 2000/20000Size� Tag  Caption
Column: 20ViewPriorityPSize� Tag  CaptionCharacter: 132 (0x56)ViewPriorityZSize� Tag  CaptionEncoding: UTF-8 XViewPriorityZSize� Tag  ViewPriorityFStretchPrioritydTag   UseSystemFont  TActionListEditorActionsImagesEditorImages	OnExecuteEditorActionsExecuteOnUpdateEditorActionsUpdateLeft�Top8 TAction
SaveActionCaption&SparaHintSpara|Spara fil
ImageIndex SecondaryShortCuts.StringsF2 ShortCutS@  TActionSaveAllAction2CaptionSpara &allaHintSpara filer i alla editorer
ImageIndexShortCutS`  TEditCutEditCutCaption	K&lipp utHint?Klipp ut|Klipper ut vald markering och flyttar det till urklipp
ImageIndexShortCutX@  	TEditCopyEditCopyCaption&KopieraHint,Kopiera|Kopierar vald markering till urklipp
ImageIndexShortCutC@  
TEditPaste	EditPasteCaptionKl&istra inHint0   Klistra in|Klistrar in innehållet från urklipp
ImageIndexSecondaryShortCuts.Strings	Shift+InsCtrl+Shift+Ins ShortCutV@  TEditSelectAllEditSelectAllCaptionM&arkera alltHint%Markera allt|Markerar hela dokumentet
ImageIndexShortCutA@  	TEditUndoEditUndoCaption   &ÅngraHint%   Ångra|Ångrar den senaste ändringen
ImageIndexShortCutZ@  TActionEditRedoCaption   &Gör omHint&   Gör om|Gör om den senaste ändringen
ImageIndexShortCutY@  TEditDelete
EditDeleteCaption&RaderaHintRadera|Raderar vald markering
ImageIndex  TActionPreferencesActionCaption   &Inställningar...Hint5   Inställningar|Visa/ändra texteditors inställningar
ImageIndex  TAction
FindActionCaption   &Sök...Hint   Sök|Sök den valda texten
ImageIndexSecondaryShortCuts.StringsF7 ShortCutF@  TActionReplaceActionCaption   &Ersätt...Hint2   Ersätt|Ersätt den valda texten med en annan text
ImageIndex	SecondaryShortCuts.StringsCtrl+F7 ShortCutH@  TActionFindNextActionCaption   Sök &nästaHint:   Sök nästa|Sök efter nästa uppkomst av den valda texten
ImageIndex
SecondaryShortCuts.StringsShift+F7 ShortCutr  TActionGoToLineActionCaption   &Gå till radnummer...Hint/   Gå till radnummer|Gå till det valda radnumret
ImageIndexSecondaryShortCuts.StringsAlt+F8 ShortCutG@  TAction
HelpActionCaption   &HjälpHint   Hjälp editor
ImageIndex  TActionReloadActionCaption	La&dda omHintLadda om|Laddar om fil
ImageIndexSecondaryShortCuts.StringsF5 ShortCutR@  TActionDefaultEncodingActionCaptionAnsiXHint$Standard|Standard systemkodning (%s)  TActionUTF8EncodingActionCaptionUTF-8HintUTF-8|UTF-8 kodning  TActionColorActionCaption   &FärgHint   Ändra färg på editor   TPngImageListEditorImages	PngImages
BackgroundclWindowName	Save filePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:09+01:00" xmp:MetadataDate="2022-09-01T11:01:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9b109123-2f71-2741-a4a3-be6c7d3c52fa" xmpMM:DocumentID="adobe:docid:photoshop:df50c30e-6172-5042-aa51-2de4f0854853" xmpMM:OriginalDocumentID="xmp.did:b11583d4-c3a4-fd4e-afca-25c912339e48"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:b11583d4-c3a4-fd4e-afca-25c912339e48" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9b109123-2f71-2741-a4a3-be6c7d3c52fa" stEvt:when="2022-09-01T11:01:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�2�  �IDATxڥ��N�P��1q�.L���w-7����(�5l�����AD@��ȭ��� &c�O��MqՄ�'sz2��?g�"� �` �+�4��'�m٫�ii�}�($��l� ��E܋����JQ�`�}� �\���v�L@����b`���U���]�d4JA���B�Q��s@QFÖCW ߍ�J ��q���&�w 1%S[^�p�F�M��]��:�i���9��o���?X���[��9#�o[�1����!��z�jhl��o_?p^��S�z���]"G�˂�E�	�	�3�J����F��1�e�h�B�lϐs(ץ���()1�Q��6|�'K&`5�DK�Ö��Åw�v�<b��h��Jh�Z���%��026'�F��؟)`+�Q�i%V� ��A,h��C    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data
x  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:12+01:00" xmp:MetadataDate="2022-09-01T11:01:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:829a5660-5e4e-2b4f-9c87-e37b8c9912bf" xmpMM:DocumentID="adobe:docid:photoshop:80ce2a0f-feb6-c94a-8ea8-39bb8ed53ea1" xmpMM:OriginalDocumentID="xmp.did:e2d3c957-f02d-1b41-8621-27da861abf2a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e2d3c957-f02d-1b41-8621-27da861abf2a" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:829a5660-5e4e-2b4f-9c87-e37b8c9912bf" stEvt:when="2022-09-01T11:01:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>P�b  UIDATxڕ�[h�Q����_݈�6*b,J�y_��� Js��ڴtl�`] ؛�S���^��n���Y��u^R��.��x�_~�����Á�9���{���	!c��7|��Mu��"�-���?ϖk+��O���\����L��LL�$�Y�����Z���n���=VCE�w��Eb�Sڞ�����E��0��a�g��7� Ca� �z�Q�9# y�w��l���;�Ɍ�5��ðM�trq��W�����Y��
$(�	)�Q��_n��Ci�N7� 2Ē�C�k���"���ui�!��`t�)h����@XfK�g��2�mtf^�$L�j%����Ъc�<}�u�d9C�W�C�9�R_���E�dV.W.b���E�Z�fX(����'�k��R�BUEx�~(�{��k� �<�H�g�q�6�@�(��
��IX�Xt��u|��^`
��Ζ��!�!��]}�̃�co��(A4���lE��I�+��n����j���_~��l��+�=�\%�E��]�2�F�xH�5Wh��7O���N��#���.���K�m��y�ȳ��`�������
�7��e��k�    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:14+01:00" xmp:MetadataDate="2022-09-01T11:01:14+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:92c47f71-a37d-f449-b661-afa4aef2bd83" xmpMM:DocumentID="adobe:docid:photoshop:1d5f6120-868f-214f-870f-25e2fd05be8b" xmpMM:OriginalDocumentID="xmp.did:ff898e28-92d8-9f42-a581-535097e6eb5c"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ff898e28-92d8-9f42-a581-535097e6eb5c" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:92c47f71-a37d-f449-b661-afa4aef2bd83" stEvt:when="2022-09-01T11:01:14+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�7~�   �IDATx�c���?��Y��3`��@A����#8 H/#̀��X�9�3���|���'.C�����}���` ��l(�����J��]4��h �8Q��J(f��P�t���JK:'!1��̴$V�����0m�\�14����b�(�� � z���J�xC    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:17+01:00" xmp:MetadataDate="2022-09-01T11:01:17+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:40a850cb-6941-0349-b059-f56f0e0b6177" xmpMM:DocumentID="adobe:docid:photoshop:de8f579b-5d7f-1f46-8e25-cfa07ff603fd" xmpMM:OriginalDocumentID="xmp.did:83ef71b6-dcc7-2240-a02a-a51d7f790ede"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:83ef71b6-dcc7-2240-a02a-a51d7f790ede" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:40a850cb-6941-0349-b059-f56f0e0b6177" stEvt:when="2022-09-01T11:01:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�   �IDATx�c���?###2��G���?c���l�ϋp �^q��Q���A$(-�%/%'��������3�=�r��[ ����z�1<�0�D�O �$h`,��ʯ��R����s�C{3���;��i�v������j`$���-
��������O;�>c�������{�+��������� �_�2��p�b��E�� ��,i�4���\W���������e(j�4���\���X��_��������_���i;��C5 D�U�n������{�����=+-�X�L�@X�|5��?b"C� �H�_fZ3X�*����P���6`W��5P]�`����Ӏ�Z$�`[	� �\�l)b|�(�l�K=\���A`�̹� � W�^��q)    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:21+01:00" xmp:MetadataDate="2022-09-01T11:01:21+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:439a39bf-ec6e-ac4a-a1ca-11ea370dcb2f" xmpMM:DocumentID="adobe:docid:photoshop:a5880379-6975-4744-b7a3-812f0e0a3c3d" xmpMM:OriginalDocumentID="xmp.did:2032e218-1ed0-3a4e-ad2d-db47cde73ffb"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:2032e218-1ed0-3a4e-ad2d-db47cde73ffb" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:439a39bf-ec6e-ac4a-a1ca-11ea370dcb2f" stEvt:when="2022-09-01T11:01:21+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�,k�  �IDATxڕ�=H#Q�g^t���q]�
b>�56��	�I6~A��R�,�@�+��Ũ��`#v� ���b��X�q�q6.&z�i������0�Dyk^�b�7�����d�$�Z�J���;����w�X�WRg�7��e�Ӆ8�U�@P�+B�����U$��6@�5z��|.A�i �[ Nr�&KV��ҩ�����#��;z��÷�_3���X�MH�i��a�p	 ������˦�7
j�E֔�N�K}&��y�	���{���?'n�a��?@j�2a���^�'�w,�	-�*��|@D(gr<�@B2��%C�O|�8_��^�.��� �N�
����w��d�P7$��zĻ�'�
�#����*d�@�OC<�)#��ۯwX���͙�x��|�,����򱗫���G�?RY�30�$r���s����P\����	!~ڀ߮��k�q�O�����h    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:24+01:00" xmp:MetadataDate="2022-09-01T11:01:24+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:3afaf7db-0640-ce4c-b6fc-15db17b69e43" xmpMM:DocumentID="adobe:docid:photoshop:efa1c113-f7e9-9f4f-97ba-3762b9146e33" xmpMM:OriginalDocumentID="xmp.did:2cbebee6-769b-894e-bd65-0e34160b535d"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:2cbebee6-769b-894e-bd65-0e34160b535d" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:3afaf7db-0640-ce4c-b6fc-15db17b69e43" stEvt:when="2022-09-01T11:01:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  uIDATxڥ��n�0��Bj�<��6K��҅��yx�NL	��@�VA��v���zN�UK\U�(���'�%��@�iй�Knp�Z=����E����6.jAt{�p�G�/t2vH,̮x���Y�<�e-�L���z �0�I��]0 ���f���:Sѝ�=�0�  ����F���s^�'�E��O7i$j�4%Z`{�LPKT$��PPI�v
�++%<��IB��o��n3�'�?��Q/�-M����]B[��M�ľ� �,=o�kT�`���y���.˾�8���)°/�Oӱ{bK;����f��q�\�)�a(<v�X0���[�ʽ�
:װ�J3w�_�n(Ѓ���l��7?�%�	����j��+    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:46+01:00" xmp:MetadataDate="2022-09-01T11:00:46+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a1cb064b-38bb-d143-aca5-917a4f08a7cc" xmpMM:DocumentID="adobe:docid:photoshop:37c98265-f6fc-1b48-998e-ab64cb46ee56" xmpMM:OriginalDocumentID="xmp.did:7460783c-7362-1449-9e0a-d4169f0168f5"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7460783c-7362-1449-9e0a-d4169f0168f5" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a1cb064b-38bb-d143-aca5-917a4f08a7cc" stEvt:when="2022-09-01T11:00:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>b%��  �IDATx�c���?%�d��Y��2%3-�n �C�f��,{��a�ӏ�?�d`��Y������	���g��������������?�����=I�pA��\yΰhH�?C��8�w���#������,��0�R��~C����۟2Ԝ{�p��Ws�E�
� ��������5�����,D�;*�7���s��>00M��f� �C�?3~�l�g%������n�-p�M0�ap�<�{̰��{K	�<����u�m��ی���|������� ���;�?� �Ƞ���p��vf&�/��2���5���}����3�z������!PI��蒊O���(�ɂ?�J�e&J  ���mG�&    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
D  �PNG

   IHDR         ��a   	pHYs  �  ��o�d  �IDATx�u��kA��l6�ݴij�&1K� ����
<�VK�"�`QĿ�@	Hz�7Uk�$�G�Ń�lk��6M�$ۦ�����gW����0�}?���y��枥n ���g��l���խ�����[����	A��g�3C��z"sL�Ă��K��d>t�3��q�p��.j W�.��H7֪@�j~i��y�	��oo�X3XjP�`��T��r!`�ib(мc$��#klc�b�b �mLM���TS�ihS��;���S��w�9!q�4X-} �^"�bs�k�$!�b,�u�4���Tg=��k�eګ���6�/�җW����Kn\
7�p�b�.�m�C��W�O-ʞc�Y��~�E�G���;0ˏ��_7�]x�����弆-L������B�L/B>��kq�Ѱ�,���bр�/�
��Ǆ�J�z�Dw�\w�a���[>�&"A�+��2�c�PV5���,%�<s�F;W�`�k��ޯ��K�
�0����\�lL���&�U9����y(/|t�uN��Ln�}Q�Ň�ꊱrw� 3� �� �����	�uX]^��qQ
p�n鄕^�a�2�g�>���N�`��<��To3!�t���A�S���B�@��4"7�ȁ�|@�¦��i~����6�bU�7�MLF�X��v`�R�?_�7$NS�ߝ]��(�19̆	CeYc�T�K�w��3L[����%.{�$��/m9�? �}�뫱�    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:27+01:00" xmp:MetadataDate="2022-09-01T11:01:27+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:dd360cab-28c5-7e46-b96f-bfc884c107d0" xmpMM:DocumentID="adobe:docid:photoshop:dedb2bae-d1d0-3e4e-8e8d-b3657d940c04" xmpMM:OriginalDocumentID="xmp.did:cc8d8e3d-e751-5441-b7ea-16b540d18ba9"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cc8d8e3d-e751-5441-b7ea-16b540d18ba9" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:dd360cab-28c5-7e46-b96f-bfc884c107d0" stEvt:when="2022-09-01T11:01:27+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�<�-   �IDATx�c���?%��8w����o�2�y�!2,�]!B�P>,���������_�~��p��% �_��_���3���G�?}�� ��>}��
7�<� 7/��?~|g�����q�
� \�8�p�4�ԙs��S��&�u1�;��@��Iܾ������)��}c�e�F�㕏�c�� J�3 ����(�    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:29+01:00" xmp:MetadataDate="2022-09-01T11:01:29+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9cb3f928-c3c1-254d-8edc-dccb1199faa6" xmpMM:DocumentID="adobe:docid:photoshop:bac5e13a-d155-274e-8591-7cf4fe76c749" xmpMM:OriginalDocumentID="xmp.did:01e6f641-8d85-4b47-ac9e-d28f2302bdfd"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:01e6f641-8d85-4b47-ac9e-d28f2302bdfd" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9cb3f928-c3c1-254d-8edc-dccb1199faa6" stEvt:when="2022-09-01T11:01:29+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>Z��  �IDATxڥ�]H�a��y��9]ї�d�R��5�6�rVB��ЅQ�E7BvӅ�M�)}��D��w��5A��"����)As{N�䕁�{��y~����9HD�?���bk!	���oՀ�R[��dp&�����j��v}.*b�|�q��ʡ HX<!@w�9���#Q�󹝣ˀ�jʡ8�P���������^Ǆ�Z^Rl�x�=.g��d������ʝ����I NEgCƟ�m[�h@�L.�z$�j�D��mw�jb�P��c�S}�@����yl^�`�ڂ@p��r���H���$�p9{�FcJ��0:�:�� �S;��[:�g�n�D�,}A(��!?�pXB��԰2��e��}�^R`w�1�	�X,;�U"�T#�8)��B���QQ�Q_U���B�Pj3���ŧ��R���P���گ�/�w(�2[����sh6�ב�x��`�o<��Vˏ�pTAq���6�m1ϼ4t
�x3�jL]��V� I�#��V)��u�A!Z�d����A�}����!E�μ9,.+ۘ D�B"� /B����R�f����E����m�X��9���zp`M��>���a�9������_������g!/�<yC���͒���ϋ�)H�3kX6�`�E�?����s��,��i�ژ���m��k=�De���D��b    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:32+01:00" xmp:MetadataDate="2022-09-01T11:01:32+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:fdbe4b88-c01f-3e4f-be23-b453305ea8f4" xmpMM:DocumentID="adobe:docid:photoshop:9b147690-5a16-7742-a6ad-57ef59cfdc3a" xmpMM:OriginalDocumentID="xmp.did:b2de2f57-6bc1-5846-8624-5f732f23c890"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:b2de2f57-6bc1-5846-8624-5f732f23c890" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:fdbe4b88-c01f-3e4f-be23-b453305ea8f4" stEvt:when="2022-09-01T11:01:32+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�.s  lIDATxڭ�MKQ��2EA���
��(ZVTd�J��������E���G�����X�d����r��ҹM��:�X�{<�B)�_����P��<���]���o��|���FǨ"ːe	בp���%�����EŤ!�E,/͗����3>9MU5������D#eA=n(p#px�ݽ}��61��pnFVykN0�U�κ!?k�	:{�oMH]X�_��.`�QÃ��r�ށ��	�=�&���`(`�s -(�s�g�G�� �D^�92ל ������W�B�9�@�J��F�#��$�4�pa�(
��~ŷX�k'}0;5(�6�X��H�7,������FuTp�j��z�����j��m{/��    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
V  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:35+01:00" xmp:MetadataDate="2022-09-01T11:01:35+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:db512fff-5fb8-be44-aad6-6fed9d771023" xmpMM:DocumentID="adobe:docid:photoshop:f8192fe8-d929-b440-ba84-3e6896156966" xmpMM:OriginalDocumentID="xmp.did:c2720227-5a49-c642-a563-140210f9d2b1"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c2720227-5a49-c642-a563-140210f9d2b1" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:db512fff-5fb8-be44-aad6-6fed9d771023" stEvt:when="2022-09-01T11:01:35+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>4O[m  3IDATx�c���?%��b�9�f�%�4F��m���~�HI�%Z���9�|cd���ۧ�e�̞� � `�9����W������?��o���103���*��?>�a�t�=?#�'�u�oĻ@�K��������۫�?�}cЕ�b�� ,�A�������g���?����Ç�lg�}ԇU�������.���/�χ��~�g�Tb��".dlE>������l��
\�3�0�O(a�������UE�F��8�������S���I� Y����n Ѻ���� o��W��&L    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:42+01:00" xmp:ModifyDate="2022-09-01T10:58:07+01:00" xmp:MetadataDate="2022-09-01T10:58:07+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a36a8ff4-7598-6245-bc72-89b62da1de64" xmpMM:DocumentID="adobe:docid:photoshop:642ae86d-c8b1-df44-9e8c-7e4b81912c1b" xmpMM:OriginalDocumentID="xmp.did:5e10e400-4a1f-644b-8a7f-b0f05b573823"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5e10e400-4a1f-644b-8a7f-b0f05b573823" stEvt:when="2022-06-27T15:58:42+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a36a8ff4-7598-6245-bc72-89b62da1de64" stEvt:when="2022-09-01T10:58:07+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>hY�&  �IDATx�eSKHTQ��ܹw�mf4���F�1�R[�P�i�"�MV�J"w-\�sH��FH.��hH�E��2s|e�����s_�t�ut�������}?��/��K��#5��1o��e
��6�_���Ovo-=J������,E�����08&���P3a��gzr�&Z.�iN.*.y��{+��V�����#���(C��&�O�`Y����1�xl�{�q��Ý�_��Z�O���<h���$�d	���Y�¥�3��d�L:��k��B
>��)CYE~U��-�Amv ���h��C�%<��,�í�|X� ���IjZU$�=Ҧe�U���^���\;8��a�qpky..�h[D��c0u��-��D���e����jX����^�%t�|*CEgU{�K�����n/�h׈q8�WD�BY�B���KV%��Q�w�%���5�t2#\ Eb�:_�� �ɸ���Ϯ��O��30������Sd!�w�mM�-���Cfn�f�ug�m���4����C�L�/�#h�X«�D���MƨE;�Ǩ(C�@�[F�F��=���ucY��ѝ$��w�$)R���h�,29����tVg�M��E��M2��N_�Fڱr�[Y�I��5�X���U]���M���+�pt.6�9���ei�T"{$��n�(��ױxn6啳�S?��_�����_�������yc����̹��E-�    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:01:55+01:00" xmp:MetadataDate="2022-09-01T11:01:55+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:872b3fa1-9f4a-4243-84ae-4cbed8e00946" xmpMM:DocumentID="adobe:docid:photoshop:8825f7e1-14c1-4345-b41f-0f7ac4d33c90" xmpMM:OriginalDocumentID="xmp.did:0cc71f64-a7c3-744d-bde6-637e1aab9d9a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:0cc71f64-a7c3-744d-bde6-637e1aab9d9a" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:872b3fa1-9f4a-4243-84ae-4cbed8e00946" stEvt:when="2022-09-01T11:01:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>bz	�  �IDATx�c���?%�d��Y�����>;=���l)܀��X����_��������� C�2�����,�p|�=v��6$+-�Nο�ɰ�V5ëo��D�����b�Ƿ�A�}H��̴$�~��a��b�0�1o��.����f8�z7��7`� `�0 $ڕ���1C��,Qo�������0�R��?�� �������&[���N#��g�>�z��5�7�, Ω�7>q�/A���lL��W��m@��o��H�0������m����b�o 33��L2��d88�}�Ű���w?�1���gX�h~�5:�<_�p��9�fn3q�(�V!�a��NC�R9+;0��e���7?q��@�0�  ���.    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:01:58+01:00" xmp:MetadataDate="2022-09-01T11:01:58+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f4fd9337-7156-3642-9aae-7f67b020e50a" xmpMM:DocumentID="adobe:docid:photoshop:b1f9e015-7b47-6542-b003-1720c5f515a0" xmpMM:OriginalDocumentID="xmp.did:f4a6d8dc-15e8-534d-8739-fb7bbc642834"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:f4a6d8dc-15e8-534d-8739-fb7bbc642834" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f4fd9337-7156-3642-9aae-7f67b020e50a" stEvt:when="2022-09-01T11:01:58+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>"j��  �IDATxڕ��K�P��M��8
>�uic��� ��P�/�j���BEB���A|�t��"NnV�t��&U| t�"���zRh[�=K����w�s9!�R �@���q�2:i(e��2�(��>`�|��n��#J�6�cDq_T�JR݈"���ĉ҃�Tn�/�#.���dP����S���6pKT�'8�/�`O�qܼlh���f-������m"�� @�ƥ�	�G
�U�cP[��9;O�El��@~��0c\B������a�r:Pd�[e�j��-�OL�J�u��*�bm'� ��}	���G����i�6���kSD[�s�mܢCPV�O-�����l
(yPr�	�� ՛����u�K5��h-�Q:G���`�P8��ଢ�.�K�������Cc���V4m�imD�?�j'.���e��>� ��-L$    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
i  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:52+01:00" xmp:MetadataDate="2022-09-01T11:07:52+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a817fbda-1162-bc4e-a37f-5d9a48a23254" xmpMM:DocumentID="adobe:docid:photoshop:13a11dbb-5d8f-fa4c-93ae-bc443faf8e58" xmpMM:OriginalDocumentID="xmp.did:ece57a46-b0b9-724b-93a2-98923844a0db"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ece57a46-b0b9-724b-93a2-98923844a0db" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a817fbda-1162-bc4e-a37f-5d9a48a23254" stEvt:when="2022-09-01T11:07:52+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>� /]  FIDATxڥлK�@���9��C��`A|5�7"B�(�Gu���ũ��(F����&��q1���K�$1�)K�s����.�{�������p���E�h�/��g�;�WC0�K�4X����[	�셩I8Q���jÁ���8�%��C���JȐ-��	���3r��cq��o���]��]SrPn��x_@`��3q*��#]�(�f@��
\ ���~΍U������3Hɶ�+q@�D�}��g�$�h�}(H1@jؔ-��� 7A��<p�~��J͎^pnS�[{c�� ��y�\/5� ֬S���B�0,pH�N��j2���	    IEND�B`�  Left(Top8  TTBXPopupMenuEditorPopupImagesEditorImagesOptionstboShowHint Left�Top�  TTBXItemUndo1ActionEditUndo  TTBXItem	TBXItem18ActionEditRedo  TTBXSeparatorItemN1  TTBXItemCut1ActionEditCut  TTBXItemCopy1ActionEditCopy  TTBXItemPaste1Action	EditPaste  TTBXItemDelete1Action
EditDelete  TTBXSeparatorItemN2  TTBXItem
SelectAll1ActionEditSelectAll  TTBXSeparatorItemN3  TTBXItemFind1Action
FindAction  TTBXItemReplace1ActionReplaceAction  TTBXItem	Findnext1ActionFindNextAction  TTBXItemGotolinenumber1ActionGoToLineAction  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem15ActionPreferencesAction   TPngImageListEditorImages120HeightWidth	PngImages
BackgroundclWindowName	Save filePngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:09+01:00" xmp:MetadataDate="2022-09-01T11:01:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:4ddaf6f8-6f7e-e849-a574-0ec0dd5e2678" xmpMM:DocumentID="adobe:docid:photoshop:4987f2e5-419b-5648-8edb-4ff4760f5ed8" xmpMM:OriginalDocumentID="xmp.did:af4eca02-06ac-774f-a5f9-ce4c812dfd69"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:af4eca02-06ac-774f-a5f9-ce4c812dfd69" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:4ddaf6f8-6f7e-e849-a574-0ec0dd5e2678" stEvt:when="2022-09-01T11:01:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�EH  �IDATxڵ�[/A�g#D$<� �;E�DHH	Ah\/��|ڪV!�Ҳ�}��lk����� ه�dvfϞ�;�=gF��J�߀#��c�`���ڱ��aU�+�`X��p��uΚ�79G gC-��x�9� 9�%�������g�Vk��S���6�Wֲŝր�Q��_��ၗSw�Y�����l��I`������DF���q@�yk�^�%�3���0���Y�ױ�A�M�m��˰��_��T�}\��h�
X�bPk�~j��FDl�%Gc��
�J%$��H�,a��!��Ի�,���q"�����u�)|l!O��O}��#U�^��a������F�P�CG���&����xZ�C�gl,�Ÿ��bP�o�7���$�M!��U�8x,�)��f�H�A�^O-U(�zn�T�B�Q��P���%_�C������N��������)�R���o���X�X�    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data
B	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:12+01:00" xmp:MetadataDate="2022-09-01T11:01:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:831875a6-3435-174c-b9bc-5fc1c73ea00d" xmpMM:DocumentID="adobe:docid:photoshop:6c9934ee-70c2-164d-93c6-d8eeacb222be" xmpMM:OriginalDocumentID="xmp.did:1e21faa8-da05-4842-bba0-9d21a4e295ca"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:1e21faa8-da05-4842-bba0-9d21a4e295ca" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:831875a6-3435-174c-b9bc-5fc1c73ea00d" stEvt:when="2022-09-01T11:01:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>ʹ8�  IDATxڥ�[H�A�������Z��CDyYtW4*�`˔�U�ZS�RB*�^{)��nO�	����ڦ�Y��A����.&H��w�9�g������|����3�� "B`���Օ�p�»@��ׯ~���)V�����o~b�����ް�㿀>�����%>~�$Qwn��'��(�jkkyT�_�C��Ǚ�@��v�eO����4GV?X���^���QT��mW�)��ؘ@	��]��f��Y���t�G����W�z�T4�+I�n ���h��i�i�����Q��Rk[)A�{Y���$�)����	�]e�ceʥ��ʲ EQ�5�l�G�v��W�S��ll�V�c�5UcJU��ٻ��aֱI�)$����8#~�������{+�$L���]]U�7�:������T��*�(��#�K��_����[,`�1�쯮�9�`��=^n�tDg�P('�~&!�ch@ �P��"�R~kN�����o��v��I@�;���9s��?�
����A�J�bs@T\�I�c���y��?m��d�(�5�eX��N���Ǹ�Z�"T��A���Q��_��4(�����u���Ѻ8a�o�����7�_ӻ.��jx"��|L�9�d�<�:;=�I��h���J0�"���?��tctgƃ�D�4vBW��p~j�tK���������_��2a�4�
w�S����:؈�Y���=4"�Z8�k����v|
����\�p��'`Rgh/�����C�H&r���Z��e��'�a��V|
t��	q�/*2~p������2    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:15+01:00" xmp:MetadataDate="2022-09-01T11:01:15+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a0a4118a-6354-af4a-b028-1763a83efb9c" xmpMM:DocumentID="adobe:docid:photoshop:8b94faf1-c342-ba48-a404-ff119ff491f0" xmpMM:OriginalDocumentID="xmp.did:5c3462f1-cb98-4d43-9dbe-062ea0654113"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5c3462f1-cb98-4d43-9dbe-062ea0654113" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a0a4118a-6354-af4a-b028-1763a83efb9c" stEvt:when="2022-09-01T11:01:15+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>[��   �IDATx�c���?��Y��3������G �Y�0Sc�*�31˗��x2�h}�=���C�PA���?Y�ɬ�ݵ@�v!6גd ]]��$)�c��$E��MRYiIG�v!1I*3-��"/����HD^f 6I�ddę�͜Kt�"��QR�B�H�4(  M ��*    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:18+01:00" xmp:MetadataDate="2022-09-01T11:01:18+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:11091a13-9d30-274b-996e-9039b54844cd" xmpMM:DocumentID="adobe:docid:photoshop:21a13a7b-5c84-dd4e-b3fa-7041fcfc95c1" xmpMM:OriginalDocumentID="xmp.did:31a8491b-997a-ff43-80aa-5a0fc2bbb376"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:31a8491b-997a-ff43-80aa-5a0fc2bbb376" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:11091a13-9d30-274b-996e-9039b54844cd" stEvt:when="2022-09-01T11:01:18+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���w  �IDATx�c���?###:��G܅�?�j ����$v��+ �Y���K�$P�>��(���L�l�Z���r?�9������X��/<������A&�o$��)����T�(����{w>b���
30���Aܵl!��/�����3��2c�`�\�P�&��� �1��9NA�@��'��_�{K@ ���0���0��j Pn �������A<���Z��G5��������j�盕�����͌/�.�j�M��)��X�31ˏ��~�f��x�Յ�޽���@?o��;�|���{VZ�����.���;��._�����a1��K��F6�_fZ3�������2n��h 8T�� D����]�`����3���N�wU���c2\��w�y�E���b���u�p�b���..�\�xH�#� �_��'�@l%6L�9�?AӠ d  �p��ZL
�    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
I  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:22+01:00" xmp:MetadataDate="2022-09-01T11:01:22+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:eb05caba-31d5-5941-b171-c11e221fab2e" xmpMM:DocumentID="adobe:docid:photoshop:33578150-59a1-3548-b5fd-b24c3c4e11d6" xmpMM:OriginalDocumentID="xmp.did:c1a0d75d-7982-cf4a-b8b4-446bf713e80e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c1a0d75d-7982-cf4a-b8b4-446bf713e80e" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:eb05caba-31d5-5941-b171-c11e221fab2e" stEvt:when="2022-09-01T11:01:22+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>2C��  &IDATx�c���?(-��Dߏ��d�BW13���.3��@套��{1��Ȋ���db`�add��������	��И��cfo`�~�*&�J��.��0�^�~A�f�a�f]4��������g��������)*��221LJ������A��6�~�� ��İ��z�ſ�����Gw�KeL�;���v7F���@pd�����˃D��|+��;�c ���h=^|�����ót�7x�Ғ�`=@	�%�v ')�9Ǆ�8��ſ݋���@���\��w�O4�0���������|��`��_A���.�q11���b��_�n��-�T\|qPy2���n��&lbT\z�����c��_�^��-���{N����<�)��q/F�a�ʎܬ���{��Y������,��` gG��|5~�b�&O����(���m[���}���/�{q&���m���K�@�y@�Bx�#Q*->��ȴ��a�O�^g;~��R�T]��	��g  ��@�X�C    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:24+01:00" xmp:MetadataDate="2022-09-01T11:01:24+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0d0a00c5-692d-544d-b746-e9532236cd28" xmpMM:DocumentID="adobe:docid:photoshop:4e2b11ca-482a-8f4a-b409-00ab27a3e27f" xmpMM:OriginalDocumentID="xmp.did:249e59a9-fef5-8041-8b45-f5d5f994690a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:249e59a9-fef5-8041-8b45-f5d5f994690a" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0d0a00c5-692d-544d-b746-e9532236cd28" stEvt:when="2022-09-01T11:01:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?><�po  �IDATxڵ��KA�%:
A�D� � �`([`Yt�ےDUlx�T,B R�(��%J˲�^��0�l]{���||ofV��b�!��RZG'WH4[M�Ż������S�����SO
y�a �Tj0�����y�=�c �s-iyZ��C�n=�+`���/�n�g�©�\T�!g1Q�5�N;����Ɨ�4��\�AQi���햿3�Ae�
�Q)a!x*M�I�RA��TF 0������(���}LǞb���~�3s��
��p0��.@4��Zj4��K��N�䵦螚J�T���O�]�|a�������XM�#?\��#�/���G_��l2����J*6�l.����(�t�����~�/�Ұy��*�},��M^/c�mۛ���[��i�<v쬋��O'�_늵��j��mH��    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:46+01:00" xmp:MetadataDate="2022-09-01T11:00:46+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6e475de9-188e-1b46-9896-52eae0273cd8" xmpMM:DocumentID="adobe:docid:photoshop:08154e42-e852-384b-bd56-9e4e94073a78" xmpMM:OriginalDocumentID="xmp.did:81e9d631-92e3-a34b-b0e0-e410f6c9dc99"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:81e9d631-92e3-a34b-b0e0-e410f6c9dc99" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6e475de9-188e-1b46-9896-52eae0273cd8" stEvt:when="2022-09-01T11:00:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Kh�  �IDATxڵ��/�Aǿ�V�J[-UI�Jh�*v�B�"A,�p�!�����Op$ĕd����-ًD��X�R�mV���o��v~�.q2�z��33���|g�g8��N����tZ��}�#�,^#�����?�0��D�<4R1*2��O��a��g�<�% &Y���6����b��q$����?*�[�a��ܘ�{h`�^�A�o�v��7��\��d�{6`��܅q��C��8q9W0���c�ҠȄ�ِZQ��İ�	`�Ī��m�*4
�#;p�V7���=yTʰ��hv�0�㠁"�C�65������g픂��L,���[�m�߅i�\}	�ret�*E�#��\�K+�B���X�j����E1_x���9���$�
����L*l�+�]�G�2��]�8=S�#�z{9���-F6ϚZ��,	$D��|E�o3A�!b������ݴM4ߩ0�Q˹�=3T�ç|yj}�jo|-i��t�?^��:�xI    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
B  �PNG

   IHDR         ��   	pHYs  �  ��o�d  �IDATxڍ�[l�dǏ?_r��4i�4i�[(];���47	�I+C<��*xお�@}��Ą`�7P���uEhE�`hb*�i�m�]	M�fIL��I����^4������~�������-��ǁ��>������gD�?�]I=��8���[S��O2>��h�tr�g�F��L���	tp;�	x5�����Ƹ𶽁�~�0��K�$����M2c�k��cWӯ��u03�O w�p�g�SY�E�
I��P��n�@$��@W$���TZ�lS�`mLq1Y�J�Db(}�\��k�����'��C���;����~��:��Zbh�rO�_�����؃��A���J�*4�E;��	 j�v��+BF�����`�Y����$�=۾c�eV����쯘vs�+�CVL�<�*�kM���������)�wߚ���h��FF�׺��~�z�b���`�C���Iո�IPE�X*`Q*�ѱ�A��܏D�s~��<}n.��G�1� B���Qt��эF#7�}� ��`(l�R�RVdEi�v��k2nt��d7yM�lrd���6�q2��&�|�-�+��`���	��jf���Vj��M�`���)�a� ���g���pa��@H_M��$�ܰ�/�#"F��>�0�L.�rC�u��(]=���x��O�[x��%2����;�^��v;l�x����� K�Ȁ�Xפ����#�7X��g�=����ݳ�e��V�AYHc�v]�V߷b^�ۊ��6q��Bv�������h׋����J�2��J0k}Q"TJyP��`�h�XXof��[�b�ڀ�����^�s'B֕�U_���zkV4�mfʗ��^�_֛�0-5��^i��Z��4�2>�k��W|�"�^�k��1H�� Bc�4���`��ގO��#A���x��y��sn���TW��48�C��<zl�Z��;��f�f�t8�e�2�,)X�_v�������Z����=[}�<]!ߗE�    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:27+01:00" xmp:MetadataDate="2022-09-01T11:01:27+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:36058a1d-ee68-674f-a89b-e63e57f035ea" xmpMM:DocumentID="adobe:docid:photoshop:11304ae6-bb34-374d-ab37-17619e400cb4" xmpMM:OriginalDocumentID="xmp.did:cd07a371-394f-7549-bbc9-29bfcb920296"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cd07a371-394f-7549-bbc9-29bfcb920296" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:36058a1d-ee68-674f-a89b-e63e57f035ea" stEvt:when="2022-09-01T11:01:27+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>Π�v   �IDATx�c���?5#Mdddsv���_]M�����o߾ex��-CdX#�&|�P�74�/*&����/�o_�2|������K�S7�ܼm�^^^�O�>A�g�O�?1�D��%�n����~An^�?�3���N߸vn !u�p�4�ԙs��S��&�u1��;�8��z�nܲ�������(ÿ��y�+�ͫ_b��7l�FPm�&  �jfi�E    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data

  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:30+01:00" xmp:MetadataDate="2022-09-01T11:01:30+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9c787553-e6db-294f-a720-6653ac8cd030" xmpMM:DocumentID="adobe:docid:photoshop:bbff4f6c-065b-794e-b2be-69c7710962f7" xmpMM:OriginalDocumentID="xmp.did:118d4b00-602a-724e-b1c1-eefd0453f251"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:118d4b00-602a-724e-b1c1-eefd0453f251" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9c787553-e6db-294f-a720-6653ac8cd030" stEvt:when="2022-09-01T11:01:30+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  �IDATx�ŕohe��'�e��d�J6����B��k]�Zg�.i��(���S(Ѫ/��@�!���ܫζ����H�dI�J�3�uŹfu�m��j��rw��;�bA�@�{��>����{�!���ދ���w cR�p��d.O �;�W�3�� *j� �7��8�N�K��W?sjz��t�Q���a���]To��a���E��4w;�xV�ֽ�z�1 P�ӎM*(#���F���	�p@�@Ƣ�E��t:z��t֊5�_T��p6��|%nD�Gsr���c�5/�X{)���A�ZIv�"���S�𳕈ܾ�����x���N�73��TYk<�+�Ht��@����g��8�/�)��OR���'e�O�����??{��{���r�PG���r{��	�Ё�R�zיA�����l<~� �ƭS�����d;���p�y�
r�^�a�/����Eε1dx�s��6�Q=4����XiJτ�:�[{�)ݿ���]����aBf�`
WfD��.�CS��x"�\��P�2� :�\��t��U�ӯ wc	#b@�r�񝷧_�X3�\�!�����kע%��[�f�����Z����`� �N�v3d_�AO��I����F[%;�l���v�#8�D�zTޯwTY��abim��:��څz�{\���ā�#s�&`#-����Ko�y���:��|���;�X���هԔ΅���sS Ͷ��4�d;��4&���>�GG;�?o)��ikԔJ\���O ��H��v\!�ON������z����a4�v����l-����hf�(�[�8\�k�����5M5d`bUS^��v��7 K^��n�֑�G�~L.^�S�t�j�!�c��zĈp;lL���!����E�to���5���ú��� Iv�%���M��a�i�zP�+���=�	ct������_SM�ב\o;��2��kM_��BY����,;�9    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:33+01:00" xmp:MetadataDate="2022-09-01T11:01:33+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:7f0df2cb-8086-e74e-b2da-c42d155408e2" xmpMM:DocumentID="adobe:docid:photoshop:74e6b954-2ced-ce49-8786-10000e0b102f" xmpMM:OriginalDocumentID="xmp.did:e8263aa7-8446-a848-90ac-8389893a4231"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e8263aa7-8446-a848-90ac-8389893a4231" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:7f0df2cb-8086-e74e-b2da-c42d155408e2" stEvt:when="2022-09-01T11:01:33+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>6|��  �IDATx�Ք�KAǿc�`Iv���%�=(�b��Y{ڪ�M� x��_ ��A����(��K�ZEKmEA��l��u�츻�@�$���o��}������!y !�qB_VikK�b1H��hT��~r;��.����
b-tC��(P�$�#?� ��#�ʧ���`Y�,gVrB����,��.l��V?���д.4-kmE`�������jΗWW�#�s�ś�gx�7bgɍ'Tx��!��t�R{\�@_��@�u�8�"����^��~��	|��
��Rk&\ЎDC"�Pȵ@�g�f��;{�X��ϭ��0��=Xk:p����K�l�Mc�l���-�Q%\�(9�vQn��D��� ��CZw[9�,�ak��i�_	�ԍ��ʉ�[�叟�(��iZ��\/U��������z�/�z�Bw�R���+�V�`�k��^]�oSl�����OAͧ���2��|@    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
{  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:36+01:00" xmp:MetadataDate="2022-09-01T11:01:36+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f4984d1e-61dc-ea45-b258-a3ab76db3d05" xmpMM:DocumentID="adobe:docid:photoshop:b2184f69-7fdf-084d-9fbf-e0078002def3" xmpMM:OriginalDocumentID="xmp.did:38e11f32-62c8-544a-8f86-ed826d4b8fa4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:38e11f32-62c8-544a-8f86-ed826d4b8fa4" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f4984d1e-61dc-ea45-b258-a3ab76db3d05" stEvt:when="2022-09-01T11:01:36+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>QޔN  XIDATx�c���?5#�D�6s.E6`50%1�,���_��@�b �zF���1�����u��_��3o�n	ί�^�x��ϟ�>���(r!�@�@i�OO�3����!�g�������P�O������c�p�#���&+3�9��<*�H��� �Ǉ��oe��b��� +�N��<%������?Û��x?�c�{9�A�{����&7D������o:b �2���Byg1�a~�c�z�ÿ&)3|����0�se���'û۟��|��@i,s�~���������i?�GQ:�������a��g�멒S�)������2
�^b `������    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
�	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:42+01:00" xmp:ModifyDate="2022-09-01T10:58:08+01:00" xmp:MetadataDate="2022-09-01T10:58:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:473e24ca-c6b1-6c4a-9246-c342e00fab9d" xmpMM:DocumentID="adobe:docid:photoshop:2f28bcc3-224b-dc4b-b030-304b5d909856" xmpMM:OriginalDocumentID="xmp.did:b09b547f-dc93-2f4e-8487-1106b539efc1"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:b09b547f-dc93-2f4e-8487-1106b539efc1" stEvt:when="2022-06-27T15:58:42+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:473e24ca-c6b1-6c4a-9246-c342e00fab9d" stEvt:when="2022-09-01T10:58:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>8w��  iIDATxڭ��kWƟ33;3��dӍ�dc�d�(iH�(H+x�-�-�P�j�Zh{S�_ �P�`A�75��(%7����l[Z��!~D1��f?�̜�wNv�ĵ�Ɓݙ9s��<��>�eRJ�ʋ@�XӇ�S�>�m��B"�&39O�\�癑����(����Qg3ӑ�tm��4�[c�� �{��K^�%��o��C�>g�?�}�s�5�_��V�N,��,S�Qw�џ[�������G�^in�}����ވ�[S�-1_oHb��V:�*~���v��{U�ꂻ�Jo��̎;k��1'����N��`ҷ��F����*$ݘ��rM�u�B�e�䇇�����n������t<��d����'E��:�;���1\xT��?g�TT�ݒ�c�tf���r��:�3�=�lrgT|r}ʜƁO��vs'n.Vp��L�WN�����<�����m�G�t���cGS��"�O�y~'{��#�s��)D]���ڲ;{wx(�����⦪��j��+m��߲��۰�}��c��s����B+&z	L�Ϭ�������&݁�/��Y���Sp���@
�����(dڮ]�E5�woD�����=\}Rj򦠍x�{r��s�NX�=�a��i��/���/���������&�S#���m���o�FW��:~�¥�E�?\j��^�_ke��N�LD̨�� l��ϼ��Ӛ�s3�M0�K!�p�U��3;i�T.�н�[q|[�:zL�����$��wE��޶���h40i�D:s���m`�r8G
_���E�Lz�LE���au�������ۈQ�buo�|Z�E���x>?�����Z�8{h�:���-в�|������_�o�Ē08    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:01:55+01:00" xmp:MetadataDate="2022-09-01T11:01:55+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:fbe6993b-2510-414f-a867-51db377472ce" xmpMM:DocumentID="adobe:docid:photoshop:6510eeab-a9bd-0a43-b303-a458c8585ea7" xmpMM:OriginalDocumentID="xmp.did:5d1f4fc9-1149-3443-a1c5-e0b80c49eac0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5d1f4fc9-1149-3443-a1c5-e0b80c49eac0" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:fbe6993b-2510-414f-a867-51db377472ce" stEvt:when="2022-09-01T11:01:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>I���  �IDATx�c���?5#����k�_�B����#0dG���Kд9�3���~�����P����`عk/�P��{��5�Ь��#D�������*7�?�?��\g$�����e�%14����[Lb���ÿ�ؘ94�<�2�%*��0,qy� h #^�ޮe��d��\��x �uo~<a8�jî�s�ev<�I����.dX}����x3�4�:�ſ��dx��.��ϗf_/`���q��g�W,bp��G	�c/�2L���"F��;�dp��c`c�$�H"�� ����W��O�2���60f���t�)��(b{��g��hC��I�dfbfH��eP�3�4#<�2<�r���/C�J=0�c�3�[!�aף�����`.�� �!����{�/�3�|4�#U�C���G��c��`"����~��v���8�D\���S�61��z�x�:.>1�$9�@V� ��`�#0�    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
R  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:01:59+01:00" xmp:MetadataDate="2022-09-01T11:01:59+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b1858f52-07ba-f44e-997c-440ce8891b03" xmpMM:DocumentID="adobe:docid:photoshop:c2388acf-0c96-3143-baca-9a46136d00e8" xmpMM:OriginalDocumentID="xmp.did:be874ab3-e682-7d41-a93f-05bac917655f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:be874ab3-e682-7d41-a93f-05bac917655f" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b1858f52-07ba-f44e-997c-440ce8891b03" stEvt:when="2022-09-01T11:01:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��C9  /IDATx�c���?0222`��U����2� �K.n����<ab��*.���e�z��1���j��S�Z�D6Pi�E���z�XTZ|q#C&v�0��������m�����3�V �g=�ss���(�&AK&&�B�}�P={|��,��^��^������c���.t��-�������FȽ
4ԁ���5N��^��x���)� ��6OK/�(������
�qf܋�gd��f�a�f=T��a����9~��*�$��"i\>K����i`1a����^���\r��vʁB����%3� `f����+�u ������&�@P�f�@��y3��̠�@��g4��X/���������8�#JK.tye�|����?Ə���Qd C�~%U�����32����(��o $�rp��*�r/��>C	���3r�l�����޿����q���6�]�fb�dj�gd|���oܽXídBKN�	0p-j���4t)�B"��IQ9���h`>%�;�A�(    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:53+01:00" xmp:MetadataDate="2022-09-01T11:07:53+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8560e4c8-ef4b-c241-9bd3-a3c46bf4a332" xmpMM:DocumentID="adobe:docid:photoshop:6ea4459c-4b2d-0b4f-9708-d4bd33da469f" xmpMM:OriginalDocumentID="xmp.did:94f62209-878b-b144-be3c-dd3036e5ce4d"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:94f62209-878b-b144-be3c-dd3036e5ce4d" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8560e4c8-ef4b-c241-9bd3-a3c46bf4a332" stEvt:when="2022-09-01T11:07:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>tXz  �IDATxڭ�KKQ��C-$(�EF7K-Ӕ��H�J�j�/�?��7�n�"�1��FEc�x-�G��h�<�9���Eep�9|�|�� �1���8�0�؃+�����
�������-q��S�q��hB���@	�Q}i�DS�� �O�H�Ĵ:�q\��S>`��܆vس�H�0%zv�2*6��j~@j.ҥ�U`3�D��Xj���Ɂ�8۷v���3@E�r�F�z���~�Ғ[f݌�g���&.�P��S���3��4{�gb��sb0d��i�[��X���X�V���W�9�6��h�V�Q?ߕj��e�,^90��	C������rxA ����>4���(p��� �g��>�����K�<�k:S���t�����=B��y�ZΔ�An���$�?U�tҳ�3%�$!����    IEND�B`�  Left(Top�   TPngImageListEditorImages144HeightWidth	PngImages
BackgroundclWindowName	Save filePngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:10+01:00" xmp:MetadataDate="2022-09-01T11:01:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e11a62c2-e08a-ee47-9da6-26bfdcd31d08" xmpMM:DocumentID="adobe:docid:photoshop:78337c52-f4d1-fa4b-94f7-4288bd3e9f4e" xmpMM:OriginalDocumentID="xmp.did:64399d63-7451-7349-95b5-98b226bdc44b"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:64399d63-7451-7349-95b5-98b226bdc44b" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e11a62c2-e08a-ee47-9da6-26bfdcd31d08" stEvt:when="2022-09-01T11:01:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>&�;�  oIDATxڵ�[OA�g �I�#�1Q)Z��\�Qox#$>�
|�~��R�h���1��nw׊!y1&&l{ܙ�3��6���33��̙33K��C`8�m�R�q�=��)='8`�c�Z%ę���l�wgZ�6�Ջ`0�5�B>����`�g�ӁFKu�V��xo�,X��,s�`@� �j�; �lɰ�&�f��K�\����. ���T5��L����53am�L0��`��;Ȱ�����)����%}g��hC� �IS�i�.���FX0d���	��j N�	��2M���.�g�RwtH�� ���!����;�����+%دsmT��eV�#����K M#e-ңgɱV�߸���K�W�7�3�0v�%�b�~�ٳmRq^�R᯴m��������!��(>B@J�fq~l�vs���m�K*q��)gLoX���ʢ.�P�ؙ�S\dL��+�"�}ř�y�œI�'}�PL8���LIuq����~���+ξ_l�܆�S�΅�/$(8��LH�;y���wy�׽m�����6�U�?��'<�O���M󮓝��,o����Տ��=THӗo���m��p��g�    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data
&
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:13+01:00" xmp:MetadataDate="2022-09-01T11:01:13+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f2fa46ce-f819-9947-be89-6ff1150dee1c" xmpMM:DocumentID="adobe:docid:photoshop:d90df69d-1d84-c343-b6da-999883ef6c05" xmpMM:OriginalDocumentID="xmp.did:57e758f2-28fc-f54e-8bd0-3a6ab6a16dc7"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:57e758f2-28fc-f54e-8bd0-3a6ab6a16dc7" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f2fa46ce-f819-9947-be89-6ff1150dee1c" stEvt:when="2022-09-01T11:01:13+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>'�T�  IDATxڵ�mLSWǟsK��
(�m�e��b�v�]�N76����fK���,�f��,K̲M�}X��(+qq�XÇ%���d����TSiភ=W���v�����?���v�!B`����q�`\S�1���t����B Ng��\�ի�3y��s����!NNJT������D}AB�*��� ���T"�!>q��j��.���øb�bb����L|�j�}j��	S���wA ���a2+�~�~9}e�V�?���E�BEQ�h4��w,�D-IF�� �tt�;���-	�8�Eʨ���4I(j׮��E ����#�^#I��(�:���DcL5We��(�rQMVD��@" t��4t;���ΣC���=E*@ht#QQQ���x0x׀.�p���ө�9ٝ�L"���ߒ1��w8Rd���R
��ݨ	�%@TTW�N?�C�sV<���1�Q��L�Bc�W���������{�����۫�w������?����\���w��g��);t�G� --�clUM�ޛ��t���
N�r�-�&#V��T3����E�xv��:g�r�~��G����s�#�4��%�� j�8\Lyb��r*�'e�������ug�!��ʻ5���ɟb%9�Kp���α���0Z��h��#�Sc)e��x��M���Y�Ӿ<t��BS�*|�ٝ/9���������������-*��S�	����謀������1b-�8A������9��C9�ܜ�����mY�wz��:0���=͆�Y̘�tgO��P�qb8�_�7����napjT9n��1��}1���^�����kb��,�y]�ٖ�L�Z�5�mYY�{��c�!��M*�+U�����^PQ�;.��(�6��b�A%q���kKdv�� ���p���o�u��]����?���y�6y��*�v)�\��7�t�as�p 6	N7�Y�Y: ��ፗ9�C�b�� q�w���u��A���w!��    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:16+01:00" xmp:MetadataDate="2022-09-01T11:01:16+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:507f19cd-d0d1-5a49-8813-17492f29cbf9" xmpMM:DocumentID="adobe:docid:photoshop:f08cdefa-c43d-b64d-a80e-433d5f53d7ea" xmpMM:OriginalDocumentID="xmp.did:e878d3be-2917-bd4a-9524-a4f45300f683"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e878d3be-2917-bd4a-9524-a4f45300f683" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:507f19cd-d0d1-5a49-8813-17492f29cbf9" stEvt:when="2022-09-01T11:01:16+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���   �IDATx�c���?��Y��3��
�ӓ�0� @f3�,HI�ũp���,,,_~���I�%$Y�����}��,!����W�I���A� �����dV�� ���0R��|D���x F^!����O=���R�
�}��W�Ғ���R�JfZ+�|�M=�F�- %��X@����##�<�0m�\�s;Y��`���m:�,  u"i�p>.    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
~  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:19+01:00" xmp:MetadataDate="2022-09-01T11:01:19+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:14906ddb-9484-2b45-8442-6644d0089f73" xmpMM:DocumentID="adobe:docid:photoshop:7ec3cd41-3792-8b4a-a193-216e6d07aa5b" xmpMM:OriginalDocumentID="xmp.did:27d77af9-aec1-3f4c-a059-bff3046cf01f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:27d77af9-aec1-3f4c-a059-bff3046cf01f" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:14906ddb-9484-2b45-8442-6644d0089f73" stEvt:when="2022-09-01T11:01:19+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>W(k0  [IDATx�c���?0222`����r-b�����̯�b���<c ��f$d��=��3�U�`d`�����<�*��%i�X��y��A]���(P�����'�mh`�G�'�� )ad�F�,,��H�8��7�?$�~<}� �������DQ,0g�T```b���^�cر�7�F�� ���O%����,x	T%��"�X��z�\�@��oq���Z �2�����h�񄱀 �1`���@�\1F1���A<��A��n_���7I�������ܺeX-8ڌj��o��eHI��i����X�����'8+=e+�G�p� n����ۃa��=?~��힓�rł��� �o+� $���k��;�|���{VZ����_��Dw!,]�����(��D�2,����iI�p֡Z���)��6-`�[�����}�>@0�X��
3���*�>�S�?��S�]�d��0�X�B�,��Ȗ=Ѥ�;��ϴ)���H2�D�u(���b�� f�]
}�������+�^�Sh��0F�?���4|0���hӡ d �e�F    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:22+01:00" xmp:MetadataDate="2022-09-01T11:01:22+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:7c65103b-d5a4-0d44-8a9a-42dcb6a587d0" xmpMM:DocumentID="adobe:docid:photoshop:48c6fe1d-6077-7b45-9cae-d7f9d0ac2549" xmpMM:OriginalDocumentID="xmp.did:54afd2f3-29f4-974a-a0d9-07b12e11dbba"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:54afd2f3-29f4-974a-a0d9-07b12e11dbba" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:7c65103b-d5a4-0d44-8a9a-42dcb6a587d0" stEvt:when="2022-09-01T11:01:22+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  �IDATxڵ��kQ�g6?���lŒ֍�A�E�(�ؓ��ЃP�C���"�n�z�xP�M������)"i�����j�1�h�l�9�THC�Mb�.;����3���c����{a��p=I� �[�Ft�f�f�m����n'5h�������V�L�����!�I�|\5�!8�{�C����h� ���!�e�"�}*�6s�Yh�E���_C�71�E���ApX�\w��P;
�=�m=��"O�}:�g��t��ۈ8�W�H����T���2��٢��{�Ϲ?+����{�bJ 0n�i]�=^�4Ie��sn-���:���U����"�w0`��(�>S����g� ��/����;z&���$L�4�� =���N�D�lM��7-�Y>�v���e�H�( }>�o��g�^X">�B�7F�
��%۔Z����<cu�uD諵�D�R]�)���R�8E�ր9�H�J� �����{2�=�)R�~^@�4�����k�Jf�iV~�@�5A�4��K�"�^�{�� ��8�zu[C��$
���W�e�o뻫g�B�I�_*t�
��`�y�ʉ��#\.�[1��/C37M���5gl�į�J�"�F+*dZ�;����<�*Y �[υ������/u'�؎����ڈ*    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
7  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:25+01:00" xmp:MetadataDate="2022-09-01T11:01:25+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5698ed50-67e6-de4e-b657-56f95fca9237" xmpMM:DocumentID="adobe:docid:photoshop:36005e92-6daa-fb40-84ad-c97bba8fbdd1" xmpMM:OriginalDocumentID="xmp.did:c0fa3677-5d97-2a49-b3ee-329a00f847ec"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c0fa3677-5d97-2a49-b3ee-329a00f847ec" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5698ed50-67e6-de4e-b657-56f95fca9237" stEvt:when="2022-09-01T11:01:25+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>!X�  IDATxڽ��N�@�w��
���"�{(�MH�܂ĥ}��x !���D��>�6R�"UR��A8��4v�q~6�RK�8���2�;k
 d��oJ)�m��d��Q����\��/A9���նbnt���s�A	Q��]]V2�Ȫ��B �����4����u��-�L�ya��t�ozBP�����s.�$����d*c<��۶�栊��3��
���,�$����x�9�~pI��D��_72�Q��"��+xG4��?��F~|� ��l1�	@�zrBC����D�� � �%2�,�� �7�Nf2��`�� �iu�nO�'�,�xu1���_�hz��֟��	~������$ς���%�6#����ޗ[����\.��5�x!lFs�?��d�q�()`��S������Sǧ�����EI�P�Ȅ5�q���۝3����E��/f�K�����cB������g�^^.J��e¼!���N�p��z��SB?��u %@��!	��'��\ձr�#����&�Y�    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:47+01:00" xmp:MetadataDate="2022-09-01T11:00:47+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8a0ab898-272e-4442-93b1-44f6837fb2be" xmpMM:DocumentID="adobe:docid:photoshop:bfe1f4b8-13f6-2740-a13d-1fcf34f5a993" xmpMM:OriginalDocumentID="xmp.did:d8dc3fe3-1bd0-fb4d-bdaa-bd4f25d9aa67"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d8dc3fe3-1bd0-fb4d-bdaa-bd4f25d9aa67" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8a0ab898-272e-4442-93b1-44f6837fb2be" stEvt:when="2022-09-01T11:00:47+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>?wn$  tIDATx�͕]H�QƟwn�u��9�V��i�
*��(04�o�݅PAw��J��*��
#!���u#	����b}l6��t_�طo�s�^&��N�ag{~�<��	�,��%0��U���w
�&�*N���@z�R9��+k4huh���	��q�A<S Vd�L��Q"�E�	g[�C�0��w��F�|~�n��ͨ�';μ�!��!��A�р:ڵ'��g�p�%���� ̚����}O�`o�������Xp	�2��K�V�Ei����t�.��j�/�T��3W��m��RT�x���X
��I��%J攞��"@}�i��e ���$��7�hKy�]�6�� ���y<��)6��F�fQ��hJI�H�J�c�x`f^�I"�Zp�Tǽ~���_��ho�:��7��]�rq�Z���0PDK�����A.�J5`���Qv��M<<ֺj��۟x5W���=����[��{��{3�5
�d ��%/����X�~��O!{��Ŀkv�h,��dvM���N4K�,f�����rVi$�c�F���;10�++��ء�D�����qz�I��Q�V��M� �n�������)�W�6R�����R լ?&����    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��o�d  vIDATxڵU[oE��y��]���q|��D����hK�*P�?��-5R��T���
$^J���H#�x@E�ĥD�EM�$N��N�^�������N�R��V�f���|��� �� �Φ���QA�����t^��C������`u:}��dߎ��@%��֒��/��	���O�t�*�X�zAՙZ(H�Fs��rb�Y6A��R�oԦu"Ě@�w��6'�Kw�� ?�z�b�"��N��V��tv ($q43"(
�7@�
��[��n R��2�Ĥ\)(�e�04Q��K�6;<�9��G�6j `PT���]�����"SșS.��_�KX�n��9U8�K�z}膘;&�R �;`�/���=sw]�7�,U沧��,^����o��'!E:��\ ��]���Бؐ.�fxȅ;��j���E�������,���)�F�s�,�ү���TF�yɮks&M!�1��}��}�ӖK�|S���ڗ���8I1�X>1:ʵ#_ۅ�%�Q:W�=d��#*$܎����z�T+����7B3j�1�m�sKPH��b�~@P�w���\CW����J��y|���qrWc�$���2�����i�������G��I<7��y7��?7���Xi���00�V*�a�&0;�r�ά]�g'��|�H��+q����T�����K�K�:�{ ��dPH@�����-��Л�%b�b1Q���6������+�N�'H�9����c�g8�-eH�֭���/�t��=�#�!Cz�Kr�I2�	a|�I�T'ɻ��T*d����a� H���e�!W�ȶ.iM�Kw_ۦ�e��1�gY�(W�f�¹'&�[�u��Qb�`��!I��"ҚP�r�0���/�[|�a��h��	(KHÖ5�{}���4{#�;p��$��6�M^�u�9��mDհ�4���g���bm&;/�2BB�hw͖w� �/�+�;'	�;��1�U�Cp�_���Q�f�{��+�,��Y��(rЎ[亓P��s(���p�l�#���_�]�	\�o��v�T���وz)��^�N�Y1������a�8@1�	9�ܗ���ө7��y�G�Е�Z34�@�����X�ˆ�y����O�|�c{��X�3� ĺ�7���    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:28+01:00" xmp:MetadataDate="2022-09-01T11:01:28+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a5503412-bf16-9a43-962b-ef9efd4627b9" xmpMM:DocumentID="adobe:docid:photoshop:0d20346d-e716-0d4a-bcc2-5e5baf07ce52" xmpMM:OriginalDocumentID="xmp.did:34c49d2f-a26a-f442-bda4-7f6adc893ac6"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:34c49d2f-a26a-f442-bda4-7f6adc893ac6" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a5503412-bf16-9a43-962b-ef9efd4627b9" stEvt:when="2022-09-01T11:01:28+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>;)מ   �IDATx�c���?-#],`dds�_�������ӧOP�����O1���4R6�k;���<�?~|g�����q�
V0�� ����G- ͂�W�����g���;�Xb���XB�zl��srq1�������_@�����W/]@���D[`ai�0}�����%�����@~?���ߨ�h��g�]�+�,,?�ʓ�@�'����?�tDH ؒ�g/�><8�q ,�JR�Z�[  pU����;�    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
_  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:31+01:00" xmp:MetadataDate="2022-09-01T11:01:31+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:56143437-f562-fa4e-8174-5c4ef7adf9b7" xmpMM:DocumentID="adobe:docid:photoshop:a5dc6965-a848-4347-9c15-b989f8bdadf0" xmpMM:OriginalDocumentID="xmp.did:38e2b191-4ae3-cf4e-86a2-33e031e69e6a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:38e2b191-4ae3-cf4e-86a2-33e031e69e6a" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:56143437-f562-fa4e-8174-5c4ef7adf9b7" stEvt:when="2022-09-01T11:01:31+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>ц�  <IDATx�͖klTU�g��G_{�R� �%�mSP"l�b��n�m�Bm�(�|�@�*"A	*�����Vw�n{�K[k��"���-�vy-���n�MT�����9g����g��E��Ozz�ex�h�}����;[�@N�{��1�y���z�����=H���-n!ӟ�|�����4ԏ��4��jkP���t.D�����hi�ثz=5  ������J6kT�R����j[R�W���.n���XX�S�˒�v3@�s����Kh�^���3�U8��}d���T��̪��̦ZZJ��Nw�;�]
*�@�����b��9�R�
����멈���/l���R}���<�2���lLQ,=�z҇��Ĺ4�S�H5F�#�?@�^_��\�)_��^e� ��Z�Dx��@�O�9m���[i�(|����� �;���;�@C��S&Fn%nXl��3����t���(�]깝$�п4H�C~]���/s���GE�m)2|#}��Q�]�r��/д,ڨ��w�П��D6E���<�$4�.v;� �y�9�B���j?D��*t�X_We�L	'��jE�W��D$���!�I(����׮UQ%I��s�@�b���yy@���:(ycQ�M���y�����L��m�i���ޣ3g��$��B=]R���_�9���;$	�1[U�s��F+�m;F�a������,	�-$]�JG��h_l��Og�����m�T5�U��a%���|��NDܸ����I�k��1��*$�h�}�����3!�l
L�J뤎� �	ڰd��b�FGP�[3�եM�[�|-�幌dK|�~Jn�`U8*�RJ�-t�;٨�v;܇�Zo�B�b�vJ��t$),��#d0� ]�|�Di���YBOu��ʬYt�Fm��h�t�G3;��;2Y'U�7�z�J�m��J�R#U���N.ݛp?0iǵN����t	0qz��!�*�d��)�9��=�a����C���znjD/��i`���e7�Y� �����	 �M�z���q=�x�d�lߒNw	]���9I�/��&��I�Ҙ�9
�@\J���#'�}�1_�A���t����,����S�<�9�Lj�>-��"���
���ci�|���v}��9��˲�P	��~9��+�C�|��v���#�Y�]7�����t��f:����&n3ʾO�QE���%��X�c��Vp�(�	M���ik0p���([����]Fk˅�{�t������o�E�2z��[��8��4}�0�g�p'�BWUSlg�(�"�j�C�q{�� �[��$&�    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
(  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:33+01:00" xmp:MetadataDate="2022-09-01T11:01:33+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:924ed129-75fa-9747-b9c9-ce10b7da16ff" xmpMM:DocumentID="adobe:docid:photoshop:be7119b6-40b5-b347-b3db-181bf42116dc" xmpMM:OriginalDocumentID="xmp.did:59040d93-a60a-6541-9aa5-8525ad193278"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:59040d93-a60a-6541-9aa5-8525ad193278" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:924ed129-75fa-9747-b9c9-ce10b7da16ff" stEvt:when="2022-09-01T11:01:33+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>*t�P  IDATx���KQƟ����:,�*�E�e��E�~���@J��m���%�7ѝ���+��W�Q얣�̙�ә����j#�
A�yy�w���p8����ȉ !�X\Za��@ӴB�@��0��Gʽ��ܺs�E��j%]�,��\u��? 8 ��ʢ�(t]��!^����	�/n�}��d��²Ll�|e)���h��7�$^M�H�����'����ae�âvu �^����Ч/��� "�}
co���J�gZ-��@�x
���M0�Np@�ӵ#�e�!���������d��V��$��<�CO
*j���s��5��y|*�{Qq�wߵ�\J��M�V���v&�a�6�0�!-��Ro�P�T����#����"�fC06kq5ڃ�����&�����%6nn!%�ϓ��9���:��	�nc�PhPц�A[s�Ǟ�S����wu�����W�AOr87S��W��ڠ~��]C�0�/�(%cm��    IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
t  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:36+01:00" xmp:MetadataDate="2022-09-01T11:01:36+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b54f9dab-bc9a-7845-b522-83ead2681c00" xmpMM:DocumentID="adobe:docid:photoshop:6499cfd5-314b-7142-ad5d-655e77e9f077" xmpMM:OriginalDocumentID="xmp.did:8248e04d-049f-1d42-995a-fe7bea727842"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8248e04d-049f-1d42-995a-fe7bea727842" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b54f9dab-bc9a-7845-b522-83ead2681c00" stEvt:when="2022-09-01T11:01:36+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>Nz_(  QIDATx�c���?-#�-�%1m�\�،ׂ��X��31,�?r{͟߿r�:j��eH!) Y���[��1~���_�g���,���o����?3����W�� ��T�@o�M�K���������g''�&�PD��o���d���O3]��Y)�������Y�Ԅ�T��ɴ@{�u� ������6m������^��a�ua�}����l�K���0�S�A����8��x5��3|���y��3�IE���}� q��?��ޏ6zH�|����������_��p��0I�Y��������<3�MY�K��)��Y@��P@�:y�[  =�D*n4QX    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
Y
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:42+01:00" xmp:ModifyDate="2022-09-01T10:58:09+01:00" xmp:MetadataDate="2022-09-01T10:58:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:827843ae-9220-6c4e-a099-c0587cf3ed90" xmpMM:DocumentID="adobe:docid:photoshop:93eac7d7-4d62-1e4d-9f84-5d8b688ac1b6" xmpMM:OriginalDocumentID="xmp.did:4afdf616-e079-1849-843a-b06e74ab6714"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:4afdf616-e079-1849-843a-b06e74ab6714" stEvt:when="2022-06-27T15:58:42+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:827843ae-9220-6c4e-a099-c0587cf3ed90" stEvt:when="2022-09-01T10:58:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>5 P  6IDATxڵUKlE�g���n��Nh�7M�J ���@UE\@N��-�n=��Z�P��PTU��H ��B�Y��Q�#�qM���!�swg�։�-r�ʻk������������E$!���󣭠*�QJ��
�\��78��%�Z��a�#���l�<��jQ�|�)(�� 7��Yv2n�+8tB��3�C{��K����&C!_�L_�ܠ���*�7~�(�%��!��s�	;�>9s�o�!��s�"����ۍ�Ti�>��İ���N�ɳ�*I��E��F�v}�Z��CM�/�ݦ��.���$���z ���v�evƝD�vI���.�S-�`��oT����^���&����g���M~��1����=Q"�va�U��\�6˨���&.�tz�#���N�_!�֎�ej�a��6Y��$d.�|��
�wN�],\�~@����,��}��xqc3	x��)H;̓�?h���"�3p-�]������^����tO����Z��.'z�f��%8��|	䑠g{����;��|�� ��<��#�><1ۼ����Y��&U`o[ ����{c*�냇�@O@�E��SW�+I��*&wa��b�"����]��^eϕ�K��P��Q"9���-�f~�����,��́�AK��4���w��َfO�S�߆���='򻓮$@�����V�o�t���>ts�&B�qN֩�hx⊿M{L5iU�ˉxW��}aH�v_�ӓ�a�@��QN����CV�f
Q.���9}����%826[w��o'�3BT��;h*��º�PR����^<x���55�\��X�A[-T���6ըޏ;8�����_H�k�%�k�08�;V[�ИP�1�\���|�#�%�����L���W&��I��)v��Z5���	���?d�NH�m8��4d^.\�r
�ue��	�Z���3��*�Z氜�$a��{k_��u�L�z��0�����%q���DFp�༓�N�^W�\��	U^ 
`�߉!!��!"�7pS�k�w��	�l��PX&    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:01:56+01:00" xmp:MetadataDate="2022-09-01T11:01:56+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0f082c5a-a45c-a147-8eff-6da0f6971f17" xmpMM:DocumentID="adobe:docid:photoshop:88b7a1b0-6eb7-a847-81c9-cc2e1635b385" xmpMM:OriginalDocumentID="xmp.did:6354b84e-9c38-e246-b965-cd5c10ebbf9f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:6354b84e-9c38-e246-b965-cd5c10ebbf9f" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0f082c5a-a45c-a147-8eff-6da0f6971f17" stEvt:when="2022-09-01T11:01:56+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>z!��  �IDATx�c���?-#]-�>k)��*v�NO>�,��`Rc�2}���l��_���l	U-���`عk/�%T� ����(�P�@�$+-��,��e�%1�e�������������7Ñ�쥢�-`$ɂ�ov2lz0����s`Kؘ94�<�2�%*��0,qyC�Ko�2|���U6��B<���U��͏'g^ma��x��t��K�{��gXs����x3�4�:\ͯ�^~������������C��G��Tj�%BQ����3�f��w�,��h��L2+;Q���H&P�P|x���M6�tb�� 122���a0�G�`�Ӆ[Lb�>K��L���d�5$��Q���כ-g}B�����ɳ�E&������i�b���_~�g8�r=��G�e��U�ɋ��G��xΰ��t��3��������A�߄�G!��Pĝ�H>�l	��d$�@ ����E�d�NB8 ^hhn ���f0\3    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02+01:00" xmp:MetadataDate="2022-09-01T11:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:588efbf8-ca72-4045-8635-753b18ea2f9d" xmpMM:DocumentID="adobe:docid:photoshop:ec44aacf-1309-0c47-a068-6505ac8a8c34" xmpMM:OriginalDocumentID="xmp.did:10b73e4e-fbef-be48-a093-e792c80f4271"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:10b73e4e-fbef-be48-a093-e792c80f4271" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:588efbf8-ca72-4045-8635-753b18ea2f9d" stEvt:when="2022-09-01T11:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>_�*�  �IDATxڵ�_HSQ��s6��H���?���ǗM#�z����JLrb{�z�B�M��A��$�!q�DF��C>BEHn�)q�ڟ�J�%�����w�E�p�e�.���s��;�w�{.a��f
�B6�=�5�~�����a�jM*�iĉ��+�S����J��?��7N��WR����2�]������0�ڹ�s�$�ٝ�$���qh�&�׃;�{2L��Ek!���>��$��O.:[|��:�u�.ߊ��a��_k75[N�ǝ��s��C�Y[�\I ���/y",Z����0>k�juO�&4�,��$�W`���RJ���i�Ʃ��V^�{�;��2�x�2��.Q�����6��1(3Tl�N�T���,!��R�d@ö#/� N�n�AA�4o�:�]��*�!���_�ߋ���_ ަf��	�zt�c���v���x�@
M/1�K.
���*~h}�-�>�T
Z(y1u�����U�Pf1�*��Y��+�Y����΃aU5�g��*�<Z�8�B
�w{\5 �F�\+!��ؚGƂ�U�Ry|���,�!<�>U\L�a�ԛ^0*�`�ʪҙ�����5�F �Q�"� �� �0�>B޳�|F�n~� s&�Sx��C��ˉ�]k���\���L��@�Q���-R2`3�7��ৃ�    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:54+01:00" xmp:MetadataDate="2022-09-01T11:07:54+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a7b3beb0-ffe0-6f40-bf5a-a6f00ef73569" xmpMM:DocumentID="adobe:docid:photoshop:35ee1429-1d84-014c-93bb-c5dd5b6e0dfc" xmpMM:OriginalDocumentID="xmp.did:dc231782-00ef-224d-aec5-7a5e3f72cd9e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:dc231782-00ef-224d-aec5-7a5e3f72cd9e" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a7b3beb0-ffe0-6f40-bf5a-a6f00ef73569" stEvt:when="2022-09-01T11:07:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��L  �IDATxڭ��J�@�O(�"*.
"h�
��EDwn����;��]�r�F7���Uk+�("m�E@PĦf���1%�r2$������8"�+��5`L{����5�8���1)*Q���x��OWH���\&H�SU ��ߕ1A&<NZJV�ȀP�Ĵw�D@��>� +B#C}p��k�e~DX��2����؅`Q�jH�J-Xڸ���*t�lU��� <}�'�S腻6򟆵`����^�|�֋�d;��M:`W����BO]*�W@O�25.�)���6])t[bچl�EtZ� ��/� �@tZ����t�����h�ΈB� %cMS�D���Ҟo��'e=Ali
�=���PSP���x��!	ɟ�Q��)�6Ë�r�%&�ND*��E֒��:��"�W<�h`ڤ��"k��-�����;v{�h$��D*DG|������ޱv���"T4� �Ix��F�    IEND�B`�  Left(Top�   TPngImageListEditorImages192Height Width 	PngImages
BackgroundclWindowName	Save filePngImage.Data
)	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:11+01:00" xmp:MetadataDate="2022-09-01T11:01:11+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6a900b0f-cf94-8f4f-8bd4-a9a2b0b1dc84" xmpMM:DocumentID="adobe:docid:photoshop:be1d9db2-c274-3144-9505-da99ada835e8" xmpMM:OriginalDocumentID="xmp.did:d7615610-6e1f-9846-8407-a6b967902d2a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d7615610-6e1f-9846-8407-a6b967902d2a" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6a900b0f-cf94-8f4f-8bd4-a9a2b0b1dc84" stEvt:when="2022-09-01T11:01:11+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�A�C  IDATx��[OA�g%�����(�$�[/�4x!AT����&&>��ෘ�`| Z)�)��n[�o�Ƈm�;����2�h��&��9gz�w�̜Y	 �V6i�良�i]��tXPa}�}�FX\R(�����\_
%}Qe�c�!3���r��z�%1@,����zG���s��~{����M�H#�� t�rzfWK(���#��C SY˶.�A ��9�I��3 �ɬ���Z��Y0��3�g &��?��e�$��h�3 �`F�k����͢>� �u 3���` ��x���X������ tE3��� �5 �9�1�3��1�Q�R=��7�F���� �^*����R+0�X*a���k>!��V��@��FKp�W
�̓b7�,bӛ��@I^F <a�vnyM�E�+m@(�ی��G�sۚ�� ���`7N�c�d��;x�~�&���Dt�R�0��4��j�d���R ��'j>O�Z�-cM�7d�&�UQA�~	?RR� פ֔�?��51��
ӏy�������2��7��	D�l���E{4���#���s:���\x�@P�I�o`�>���/ګP�t���Jf����-�s\Q�"=�ٞ��}e[�uN����,���ҷ;��԰6��u��5f�Y�N�9�{�e���5@�$�6�ֺ!�����@�+�O��P�t��{��t+w6��m$1L@2#�N{��:�>�Joz5��׊�gP���/؊���Ո�d��    IEND�B`� 
BackgroundclWindowNameCutPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:14+01:00" xmp:MetadataDate="2022-09-01T11:01:14+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6374dd95-1033-0b48-b08c-8a8b623ecb1d" xmpMM:DocumentID="adobe:docid:photoshop:66dad3e9-784f-b244-a3be-a8a12609de3f" xmpMM:OriginalDocumentID="xmp.did:5dd6aa92-7f80-3f46-b5dc-cf87557ae015"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5dd6aa92-7f80-3f46-b5dc-cf87557ae015" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6374dd95-1033-0b48-b08c-8a8b623ecb1d" stEvt:when="2022-09-01T11:01:14+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>s��  �IDATx�ŗ{L�W�ϯ-P
>q��N�PJK�`�){D�m����2�tN�,�-K�Ð,����ئs�lЖR��a���,n>��Rp��s��b������ܖ.@P�Vw�?~���=�{�9��cx�Y,�H�2�v���I�z��@l�>�~�Zy� E�L��}�: �����+�I)e����BJ���X���a-*��aƴ�����r���hx���(b��*�	rqKiYY��PVq���
cǌ��3_R����j�\>_E��f-�4�������F���
!�l`�&H���n:�lθ�k�`4�+����E��)�؟W*ÎPBT�s|�/W3�-�-�.���k��iX����!a_�z<r"I^m|����������췉h���!
�^�!�/?�[�P�u�� !���#���c<����>+��[�*���r��n����9�m2�Wf���PTj������^a�\�	�V̔�����.h ߖ��R����^������'\'j�3��lw_ �Î(H�ƟۯC�,i`�����@�x|> '��u��9��=��;9�)"6̌҉�S��Ɨ]�����bk�-,4,�������}���t1�qC^^�"wW��u����t�'�?'�[�sg0
�$�b9i��q��[�rW��^���&���ݶ� �:�߿��HF�_�H�6.T�{'���R�G1�,\�|�T���d2ּ���Ѷm2��e��u�eMF���a����*�� �L�}��L���TF@���f���Z3�l��蔴������|
���Py���F���.
�x��<'���j�E^~�4-H(l_ְ��/�|ܞvFE����K�Ѝ> o����C��2������n����Q�t�Ś��q�z�C1	O�H4��I1�h�N4��w��J*�5��I�y+��i��� 4�νx^�ƕlu4�o���8&�?dLX��2�[���Umoͺ���GZwb��#�A����?����+��=�L훁t$"��U�� �"Sc�a���>:�j��JL�F��-:i���?ob�~WEJ�x5�g���=xN��1��S�1�q�n�~VIT��oS���+�����FL��y�K��M.k��N&jd���Y𷧋�G�!�\���r�$nށ �bv4-м? ���:����J}�}ڴ5�� a�0J��4� �k܃��!l�yӣ��y	�Wb�v�k��{����(�g�y���� X�FS�pd��މV$_��JOĄP��^�S��\LA�i��<��t?|:I�2h6*ʎ0U��5M� �~rd�Xֽ�W=T���x������6����0:�!�`$(jUxzno��:�c��C�_�_�˫21    IEND�B`� 
BackgroundclWindowNameCopyPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:16+01:00" xmp:MetadataDate="2022-09-01T11:01:16+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8dcc3872-1c63-0547-b01b-0bd4c714160c" xmpMM:DocumentID="adobe:docid:photoshop:63ac9a14-4744-f146-8a0c-f85702de9a25" xmpMM:OriginalDocumentID="xmp.did:61d9e7e8-9e4d-5142-b495-d81e8d3e2148"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:61d9e7e8-9e4d-5142-b495-d81e8d3e2148" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8dcc3872-1c63-0547-b01b-0bd4c714160c" stEvt:when="2022-09-01T11:01:16+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�ڲH   �IDATx�c���?�@FdL�5���*v�NO>B���vb8 %1�(C��_��������?��:�j���`ؾsɎ��@j_�zM�#��  �D9 d. R�C�OVz2+]B W� �H��"Tw��
< kaEQ �~bB[aE�\@��Vtl�]C [a�����B���*3-	^X�4py � xV�Y�r4�b@� �7TFF��ô�s)�������0�m;�t�@  �����?/    IEND�B`� 
BackgroundclWindowNamePastePngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:20+01:00" xmp:MetadataDate="2022-09-01T11:01:20+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8d7fe85a-02de-8b4c-8bf3-b7d3af7d8607" xmpMM:DocumentID="adobe:docid:photoshop:cba686f2-47e9-6441-9fda-e471ca02127e" xmpMM:OriginalDocumentID="xmp.did:1cfce908-e401-534e-9d7f-e49f0a6880e6"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:1cfce908-e401-534e-9d7f-e49f0a6880e6" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8d7fe85a-02de-8b4c-8bf3-b7d3af7d8607" stEvt:when="2022-09-01T11:01:20+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�!�  zIDATx�c���?0222�WW1��H5312D�����_x���F�0�_$ ;Iq���R�@%(�1��`w}^I��#���F	���X��:u<cu}&MS��*��������"�ג����L,G�������{���[9�D�' ŋ���L�(�����M����j��u�l��*6��@&@�p��ӭ��?c�H�03�C3#�����{�Fu ��Q� ���9qQ r�� B�h�v2 џ�)��W���  �� ����؄Թw�㭄pUj.qAL��$�t14�&��Z\\�&=�!%1�(̙������Ͽ,����G:�h3a\�!����w�����O�#p:�H~��M9� R���kG�t��F��%O�@ �YiIG�:�P���� Y���������Ċ��	;��"�!�+T���
��p�E�]%�B [�t��Z���L��WC��Uh{�	;��*C`Oa<T�a�$�G�4�]����A��YN�O4i;��O�h�K	;��6C`k1j���C`Ka�Хal.`<l�Y�K�/�h� B}C�6s��� �  ��߃��:    IEND�B`� 
BackgroundclWindowNameUndo - internal editorPngImage.Data
�	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:23+01:00" xmp:MetadataDate="2022-09-01T11:01:23+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:48fff082-97e4-4b42-8b5e-21b3a6e07d30" xmpMM:DocumentID="adobe:docid:photoshop:52765835-7494-4b47-a63e-2a7bfe60767e" xmpMM:OriginalDocumentID="xmp.did:a2e9940f-108a-074f-a00c-6f94f50bf75c"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:a2e9940f-108a-074f-a00c-6f94f50bf75c" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:48fff082-97e4-4b42-8b5e-21b3a6e07d30" stEvt:when="2022-09-01T11:01:23+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�r�v  _IDATx�ŖHSQ��}9�K'�P�{sde����?��鏰��to!D�a$i�?����_P6soTH����� P��Y�A8�,�m�v���kL7�ۺ0�����sϹ��`B��'`:D�8@�z�79���m����8x�V�u�R�kz�k��ق�����P[`i5� 3L�H��[1&;@X)��`�Z �j��"�N�u:�l %�j�E&��#,`2yY�-m �s5�ц�f"`"�
�ab(@�/Σ���K�>�	��@�`6S���]?.I/��̻�-�l��Xqݾd��7�A|ᦗ�6��=�ǔ�=�z�	�?F_��/s����v����>�~~x|%i��6) L��sVb�����D�N��Ơ��y��G��� ��γ�s�ǆ����]QxR�ӾX�X���G3�|<� 9g�{��c�aw��6��%����^�I�2 ��TCy�Ư�9�g�B )�CY� m�)ŋ���/L�`����M��H�~�7U��� n� (��A�����Y��(L��'~|_���a2; f{�Q}�(�"6!W���lt� 5�8Q�Dsr��ϒ���YX��ܨ��;�R��o��_�=�(��{�� ����Wo��#s Pw�F�f{ĕ�)ԏ���R�� D��N鿦��Q�Q�0�U~��
�����D����sMY7xWK��q�Wd�-o��\�3�X1u𞞓�!� tW�NL�<�u:b��^��%x� 4縀�:�ci���J��t���M��p�"��Qۗ�x� j�U!l�i�θ6Yg,+@x�V�1
	�����\�-U���6!�(]    IEND�B`� 
BackgroundclWindowNameDelete - internal editorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:26+01:00" xmp:MetadataDate="2022-09-01T11:01:26+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:36b6ce81-33a5-fd43-b16a-6538262a8fcb" xmpMM:DocumentID="adobe:docid:photoshop:a74ed8a2-6a9c-6a45-b72c-a2d3a3ac3d54" xmpMM:OriginalDocumentID="xmp.did:6815661b-3868-f949-a18c-8f9656449dcb"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:6815661b-3868-f949-a18c-8f9656449dcb" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:36b6ce81-33a5-fd43-b16a-6538262a8fcb" stEvt:when="2022-09-01T11:01:26+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>Z��  �IDATx��]n�@�w܄��TQ��@�,��`iQ���SX�#���J�V�4�!(���p��̬w�������D�������ءBr�A �PJ�������~,Bdmm����ѹ>��y��}߃�-.8��M���K�@gw����	�ķ�W�B����2<�;��q?�q�U��!�ZW򔂸)�:B@��be<�2Ou���t-jy"(8��A��Å���Y�Y�<B���p�gր� 2���"���xn 	�l���K'0!A'"v|8�ˈ�hw�.��!H��7����xa��q��	��`v�#�e��� 0Z�L��Q5���Ib���4O�VՄ��7�h�|�tPQT�ං#r:�o����t�����>��`�`��)H_jr|�16wB�k�Ǣ��M'���|�i2v����#��6Z�Y8��oDE:B����u����⭸h{Ũ�upB('�9���i��QqU�v�N;�kB`a"D�};6O j��b'�2�Nv1�H^�~��%�M�uT���0�����D+?g��G�ƫ��n��_BT](C��K��\���3k�E�Ճ_o���X�T��
�C�xf�כ�A0\����˵_��T��G< �Ӛ���"�    IEND�B`� 
BackgroundclWindowNameSelect all log entriesPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59+01:00" xmp:ModifyDate="2022-09-01T11:00:48+01:00" xmp:MetadataDate="2022-09-01T11:00:48+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:511b869f-52f9-344f-ba4c-a637b1ad66f2" xmpMM:DocumentID="adobe:docid:photoshop:deddd1a5-dfda-7742-97c1-5094c07dbbf0" xmpMM:OriginalDocumentID="xmp.did:bc5e0618-0e49-9245-9876-d10c035fda57"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:bc5e0618-0e49-9245-9876-d10c035fda57" stEvt:when="2022-06-27T15:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:511b869f-52f9-344f-ba4c-a637b1ad66f2" stEvt:when="2022-09-01T11:00:48+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  �IDATx���KSqǿg�M77���Y�i�]0�%],1F��uyt!��2{���B��B�2�nЋ��$��f�ZZkk�1w��r���;�	�|�/�3��������y6��8,��@:��k7���#��y�bV͉G���z��w�`�b2�C
��<�)e0T��W�C���s�݋dx����5��ӗ(p�i�yz W�=��ejA��Y�~��"�o���!i��҆p<!ieyhӪ�X"��`O>�I\
JB^���2	�9�=r��S0�ɥ��u%Ti)~=�ǡ�� ��P���y�p�l_k
�h�ΊY���p,!d����Z%����ṓŹ�ND@��;�`���&Of�!p�iE��@�*l��G����ꆍ p	N0�˜����Q �WO���)�d���K8�|���0���FbB[��?y��!27T�I�k�/U$[�W�}��tLuK_%���6�xC���jz6�f�p{a2R�Q���������*��T��?�$��m�4�"M�YS��M�998��q�h5��_a"m��v^jK��da�̀�]���2��������:X�x5�Gۉ�x)�h�pF��iѵ�<s ^gM�}v�i�0���]C���V�����7�����8�
�h)/����P�4ӤP{����n��J*�@K9���>�yC9��"5������    IEND�B`� 
BackgroundclWindowNameDisplay preferences windowPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��o�d  �IDATx��W[l�U?��_�^�u]�v�n��MA�(b��aLypgF�
�|VCLx����(!�D�'E�Q� �`r�}m�vk׵�w9����n�$O���|'��;���v ���/	�4���ɳ� �3�v�s䳻B`�릴��y�du�	0�`�����w��Б@+�з�3v��6pT	K��K��wV����$�zO�F^_��;2\�{�Gل8H���2����n$Y ,SJ��u��$A���ks���>�(�NAr��:3yZ�}H�,I_a�7PF0����������:l���#��ȟ"�]um���H���է�Lj�N�5����������K*��k�H, 0kb[o�m�]�U�� ��A��ߋs�J5�.��$�+3����r, 0|4���~m�� �/ Z��>����H_��T�3�ײ�r�ܸ�x�wp
��q������c�����á&K�t%�@�U8a8���/Gr�Θ^kJ��%iw�!��!/gD��k��Ϭ^������6"l��a}��TsC����gӜ�o��Y�������H�!B���V[���� ���<5ؖ����<h�6�>��a�;ЎKo�;��T+�=R�x�K���J�:�i	>'Ev*I3��	J��֮�PEǛ^���V��z69�jSы��ĵ3��W�c�X���v��S*�(Q�T*��u�t��ޖ��2C������Bz��p��D5���+��Rz�%l=��7�*9*1t����;Ƭ����Ƈw-���Ӳ	����Dv)�����Z9jh�V�S�h|p!����Ѿ�o�@}����Mh	�5[eIvT��ȵ����Q�Ȗ��R�Ni�P��#?�$Y�>�������W�ө�9���|������ �զu����r��',Cd�|�]���F��E����O3J�\*Ɵ(u�jh�湜F39�$���p��@�0,?(�K�s�U[�x!�����5�G�r��S�"�k9�k���:�p[��ځ��4��	]e�?1�,J`6�+J�&kiU3ӫ�٦S�c�l2F}�~�Є��\.{��泩��x��5=�fũX�\g�5�;�����Rzx�8/�>Q9���<�(�|12�/I�Y������f-1G<����˱ِ�{���E.�j���e�E�B)@�s�$3`�R�|Cb���[����}6I�D=���t��0�N��j�W	�A8�:P���P�q��v�6�g��*��Z�r�³E��/0U�2�"ޓ�֭������|N������ܤ�	!X/� �8�ZSZ$!�r���e��o�	�\RꪫJ5�%5�PyY[>p4�b ��5޿��=L�7��5vƼ�^�S4��1vg&���e�x���sK�Ȗ�i�;O�;9�9�d�:]zj�    IEND�B`� 
BackgroundclWindowNameFind text - internal editorPngImage.Data
v  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:29+01:00" xmp:MetadataDate="2022-09-01T11:01:29+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e43091c6-e8cb-0045-bd75-6a24aa23a6df" xmpMM:DocumentID="adobe:docid:photoshop:a9c1969c-261f-6249-b22c-7941c9cab274" xmpMM:OriginalDocumentID="xmp.did:ae86bdf9-ff55-d54d-800c-03f6e672ba6b"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ae86bdf9-ff55-d54d-800c-03f6e672ba6b" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e43091c6-e8cb-0045-bd75-6a24aa23a6df" stEvt:when="2022-09-01T11:01:29+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>n�F  SIDATx�c���?�@�A� FFF���m;����0���2|��	�?3|���!&"��C�5l7�t���2p��2�����p�Ƶ+D9 �?��w3F0� �۸忐���� ???���ߑ0�0~\tV��j�4�u�srq3p1'ÿ�~��Ŀ� 1�·�_�� R� ��V��b�b���e���+��/_��h ���Ë��i뀹3�2L�2�!?'���������!���aʄ����Q�:`��Тx�+�Q��k�-PF��ܒafaa��Ԃ�	�B�SP��O�X<Z�h͆�$�Έ�H
���:  V 6ޣ]    IEND�B`� 
BackgroundclWindowNameReplace textPngImage.Data
E  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:32+01:00" xmp:MetadataDate="2022-09-01T11:01:32+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:fea976a6-d234-7344-8c9e-dc0b91c0773d" xmpMM:DocumentID="adobe:docid:photoshop:ff312be5-1fa8-8640-aa5d-0b62de7111d8" xmpMM:OriginalDocumentID="xmp.did:ef1bfb0b-9096-ec4e-b88e-3ae35c43be82"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ef1bfb0b-9096-ec4e-b88e-3ae35c43be82" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:fea976a6-d234-7344-8c9e-dc0b91c0773d" stEvt:when="2022-09-01T11:01:32+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��[�  "IDATx��W{PTU�ιwaQvA��2���j�(� �@S�eӔZV�f��=l��ǌ3��-+��va�g"�f�C*|�d>�p�Ų��~�.V�F˩:�e�~�;��;�{]����{�1zUj��_�Zs���� .F������BR�у����	��Ԭ��c456l8�e˖�?���3]��.��x�|����& rq6^?�3I�_��|w�����{?#�D}	a����8w0I���$����A �F� �b)� m*���1������1Ne��=�o������zє���"`����V�}$I.�{\�������S�$��^�KKK����=���E�H��Pi+U${�x�G;7%������|i��%F+�?B� (l ������\8���k/@�Pౕ��TX�h��I�2OO��M&��CI����,���	�����Y���qyN��۹����p���G���PAz��,XS���^�0�8���'�� t%���@Sh����}Ne�f�ooxn@�϶	_G�ʉ��$�����A��֥!
Ul�z���zJ��R���H�P��v g�xƸ[H��z�ka �����ˤH)�x7���Lg�8X��X�󖗴'�b����N�B��W�7�p��n0&?Y=�aD�� ���qe����L���p�������4<�xJ ��ü9R�\����h�`�}/׃K2*^3&��9����B�q37|�|(F�1r`{Ib�߃" 쁲x�Y��8[%\����U}~ֱ7u����2����)�C�_L��YY�U���+�*uD��iߢ��v��'dӄ8RG�|PH{�Y�!z�E�j
���|�/���
6�zq�j� dh������b�+��|�~[���_p�7�k��@7B�.��
�c�
����fC0kDh�ʑ�[�UTm��64��f�ٟL�����5��T�8��_�~��=%5�R�t��)�,�����X+ �I�>��Fbr�ʔ�Y}kl?�*50)�ˇ2ŉ�_e2ȱ�j�p�q�0)s��)|6䢝�xC!�Z�3��A_Q}�V�40-j�:h��I���X�ecscڽ|؉(*z�(A6�CZͥb3Z�t\B�������jS����v�w�F�IL�"E7�ަ�*o�L��A�w�F���+�O�m P� �w���a��s,;�T�#M���;\��%�²=�i ܳ�a�h�M$;jZ�6E�B`��M-�����$�=k�)\�'c&�E��2-��$!��n=z����JWm��3�9�>W�`=�R��v���h&nZ�����M�>ȸެ��[ �GQք�P�dF*�*��d칬[6$`�dz�T�q�(��+%�3@�'�@����&IK�SE��yD������n����	3�t �]ҝ9E�ʂ��P�ҝ Qo�h@*\�B
i=�Ҿ�0��z-W��C�����tr�"���;<#u��_�*��3���*��H�.HU�����O5�T�9��]�S�*:���Ԛţk��C�[��Q�g��vO!��C^rn�b�c��.�3��y�����둼ߧ(��Va��ϊ?����V��������9˘�����1����	����ԤP7��^����bP�/�y����ϱ�"ɨ��N�<�u8���x��%g�`�i�L8T�6�B�@~HZ�HF&�����c�-�lD�>�R�c���z�ȃ��`�`�'.���}�m�F<!(ޅ.��_Q�nFvއ���<�M��FP��t(@D�n�^(3S�Q^,�K��s  P�H���=�    IEND�B`� 
BackgroundclWindowName	Find nextPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:34+01:00" xmp:MetadataDate="2022-09-01T11:01:34+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:16e01967-c303-f546-8650-184397ea53ec" xmpMM:DocumentID="adobe:docid:photoshop:f739d9d1-ab02-5641-9911-8f1f05ce751c" xmpMM:OriginalDocumentID="xmp.did:23eebcfb-a089-9d47-b172-cf28c2ad2c51"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:23eebcfb-a089-9d47-b172-cf28c2ad2c51" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:16e01967-c303-f546-8650-184397ea53ec" stEvt:when="2022-09-01T11:01:34+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>kjd  �IDATx���KQƟ���~��Κ�d�UEV��XTta�ua!�B�EAI�T$��EWQATP�kR���E��L�sNgV]�v�uc� ^�3������w�CcX·� ���Fo� ��b�$i>f!�J8��L�]�F@����
@�T蚖�#ÃE��xV�4V V � �z�X8�(��BPUuQ�A,�mm)R�F`��-��������R
�4x�H�XX�1*P�ƒ��؉h4�h$
�ZP��@�3Y��%�(/�����}��N���K��8��3��z͇��� �:�z\�ǿ< ��W�J^X��A5ay <
-Q��F����x�,�<�
��uP߆� .�3q�N����a:���s�33����Ɂ(t��Pw|��� ���LP>
��W%AJ�Zo��"vd,�3��y ��1�?��xċ����kK���v��o���ؙ�s�|.�����C95, � ξ�&G,�7��ƃ���r�<Ǧ��"��8&Ucj�2w
�r'c;��`0�d��n;�g}�N�gM��;��+�s�7�qep. ��>W��س�A����5��f�0�@�Bĵ{c@ڝ�Q6 K%���h�;��h+��j��}v]�a޺��~~�<8��]}Y ��řJ��ۧ'�T_��d�=b��� ht�y���     IEND�B`� 
BackgroundclWindowNameGo to line numberPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:06+01:00" xmp:ModifyDate="2022-09-01T11:01:37+01:00" xmp:MetadataDate="2022-09-01T11:01:37+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:aab97ea8-bb47-c04e-924a-0e3708646566" xmpMM:DocumentID="adobe:docid:photoshop:b2cefb4d-cede-fc42-b244-d702032500fd" xmpMM:OriginalDocumentID="xmp.did:92d6509d-d45e-0c46-b1d8-d0555401cfa4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:92d6509d-d45e-0c46-b1d8-d0555401cfa4" stEvt:when="2022-06-27T15:59:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:aab97ea8-bb47-c04e-924a-0e3708646566" stEvt:when="2022-09-01T11:01:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�^�g  �IDATx�c���?�@�Q��U8m�\���$�$�R��9�Q�[���߿d[������8HB@���5��~˺��j@`p�����?���/�bb@�(�? r���@�x7��_�W�u�-�������`NL_���Wy���ipo���{n��[	Hh����0ßԛ��7i��o��?,@����@�x�ʫ�i��~�$tvހ��`@v�0}.�����`�;@{���0�P-�;$��un�j���x���K�Ŋ��0003C������G������B��+��4�-��#|���~ �[��|�A�4��	� t���s����'ݏ�q.��x)��7 ]~��:������������z?��!�b�9@m�P|���_��p����,
T�\^�����af/�iT�w��j)P�v(��шw  ���W5��    IEND�B`� 
BackgroundclWindowNameOpen online documentationPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:42+01:00" xmp:ModifyDate="2022-09-01T10:58:10+01:00" xmp:MetadataDate="2022-09-01T10:58:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:87dd2bba-2fa4-6141-8eac-e2fe8e15c9d5" xmpMM:DocumentID="adobe:docid:photoshop:c7208901-8e88-a14c-a5a7-593309584f83" xmpMM:OriginalDocumentID="xmp.did:47a18cb1-f8b7-1c4b-9d99-4a76f1c61a69"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:47a18cb1-f8b7-1c4b-9d99-4a76f1c61a69" stEvt:when="2022-06-27T15:58:42+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:87dd2bba-2fa4-6141-8eac-e2fe8e15c9d5" stEvt:when="2022-09-01T10:58:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>)JU�  �IDATx�ŗYl�U�Ͻ�-�t�ЅR���%iKߐ��$`� �Bd�L (�cP�X��@P�Hp	ЊBm;�"J�R��tf��z�e�3�3�Y������sϹCc�(/� �$�e�)��8k>��b��q��y�9J� X708�9��v��[*%3i��	�6\ʠ<�L]GEB7�Ɖ(G�p� Ma����
�2�J��=L���\Uy���%��#��l^�q��QcC��i�4
���}9�bdM��Ε�L@]-.yn��W=N�M$$9�3�U�A�N8�4���v���%��K���D��'
Vnk*��5Y;�"ƊH(��P�.����B��$��ET��87,��8(���zp�{�oP��qzH�BO`���UWlU����e6�4d��V�#p�{Z�:��9P5x��-8���!�+���;R=��sEŗ#�.���]�D1�W�T^ ^;�W4i�!,r�p��~�@��-G��+�c8
��'��`�N1�ݕ+��b�zb&�6)�t>��݆��}����S�.5�O��MWn��#�"�+�f�j�7	�v��R�}��u��m5�u��GgB��\�w=��jw\­��	���zN�;�1n䃪oQe��v-�m]"�����g�ӕ����]vj���p�^0
��`�v��5��?���G���AUf��kʿ5L9|e�3�_#f�	���{���f�a��x=�?v�ȅE�fe�J��'B�~��@j������niM�w��%6� 0�%ƃ�|�5`nv�cD6�G�=p�w'!�Y�[(m/���8�җ�u�)��gc �aY>p��~���] �ZB����~�����c
hja�S\1��c�gg�����QxwH�/t���<*<f7 
 QX|�Dw�x��[���X	����!�:ݑ�W�`�͖��L̀��M�V��r&h*p�]���v�ﭮ��hJp��9P��n|�����n�gq��p�*!56	���ˢ�K	��옙���m�����BO`���|��ت�F_u�J+�R��UZ��9|h�4X�+��a�^R��<��?�!5�-riGu�	��K����$�e��v�܈?
�fDK�ٌ.�ϻ���L^H��xl�J�vl<gn$���$M�T��_3�͸nX��|��pu9���(IW��SS!G4���|�~�M�(<ZR-���j@
o���;�@R�ty��3�8�tl�����WRC��W�ճ#5g䑬�����Z;������ey�Ԗ��p�{�)hX~(��V܀���֨�Ң���6�>���A"�1A��tǭ\Rà�9_��yI�1"v�p����#G�F�;�o�zCj����ؼ��a�9��\�jx��lga$���|���_3lw[(%��+l���1Q�nG/��w��Jx�=�G�������%����� �X�ۜ$��Z7Z:�9��N��?�6!����    IEND�B`� 
BackgroundclWindowNameReload filePngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:01:57+01:00" xmp:MetadataDate="2022-09-01T11:01:57+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5ee772e3-fe24-6347-a76a-2672227d635c" xmpMM:DocumentID="adobe:docid:photoshop:aab72e79-7ea8-1147-b968-3b4c65c1432f" xmpMM:OriginalDocumentID="xmp.did:23708d60-cf6f-b642-9b6c-8fce8ef2b3f5"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:23708d60-cf6f-b642-9b6c-8fce8ef2b3f5" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5ee772e3-fe24-6347-a76a-2672227d635c" stEvt:when="2022-09-01T11:01:57+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��c5  �IDATx�c���?�@�A���Q⢿@����G�Ib�,V�$ƒe����XXX������#�� _o��;�`u] ����k����@ �#�� l���������0�� <�OfZ+M@�q@0R�w?�1{�����S��|b`g�bP��c��b��V�9�|��G�Z��S���fXq�	h�,���2�K2�	2�������`5֒!	�k�-qyC�,�:�p��!�O�
dy�PBeӃ	{�����þ���瀹��?]�����)��3zο��0�R� �8ÛO����n3��b��gHך���=O�1��F��O�n�?fS���40l{8�a��ai��=��p��q�8����?_fW�c�P-�:���v���9���7���#�a�<�.J)���x�PpĐ�_��!T��z��dP�3�%�U�b�:`��pQ�my�A�K�:�a���%C��Cw�Aʮ�n�3�˥3Ī���Q� '�8�[O1<�z��Y&\�K��<�r�aݽn�ӯ63�	;1,e`fd�����B�+�(e8�|X\�S��������o<c`bd�a*5�S���n.2I��`>(��X����%��0p�0�
�1XK��kH\`d�;��CQ�7p  ��/�G'�v    IEND�B`� 
BackgroundclWindowNameRedoPngImage.Data
|	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02+01:00" xmp:MetadataDate="2022-09-01T11:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:2b3b1bcf-41ba-f84f-92f1-79cf5f93d248" xmpMM:DocumentID="adobe:docid:photoshop:8a03faa9-25f5-5241-b953-9d294ff0f551" xmpMM:OriginalDocumentID="xmp.did:d050376b-8c71-154f-9441-600a82ef4849"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d050376b-8c71-154f-9441-600a82ef4849" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:2b3b1bcf-41ba-f84f-92f1-79cf5f93d248" stEvt:when="2022-09-01T11:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>:�?�  bIDATx�Ŗ]HTA�g��(idKA��j�C���>K�H`D��?�EE��YD$�����a�!$,�|�o�K�۽����P�[w:w��m�n�ռ�0sg�oΜ�s0!�O�� �j@��� *l�A��U'eȥ7h4��!֬/����_Ia�	�p	�D�E��L:�����H������f=�����Ы�oQ"c?��E���@� �jN�ՠ�#�O��V�l� 8Z��^�wN���S|����j���JFGaN�o̃�>��ʼ t�������i|��I��Y�vt)�yK���ˠ9#�w8��
9�t��nen�f,��xg�?����M�+�*�>�������5AI ��A=V(Q�(g1�J*�j]Aa="���VI ��g�Q��}�Z;��w2W���K��)�(�*n���*� ���GI�kq�@
E�}��Y���E��J����,����
)�jX쾇#Ȟ�t�0�ꙤoD�4�C?�`k��6zNVC�F��ֹ ����]3 �k3^���x/�'x�����Z��\ŵ�,�Օ�x��
���֢G��s27�?�׿9L?dȼݿ,5MŅ��#|>:�,8� Z�s�B�V	y����B6 !�Ab�J*q�;����[�|� $�9���J7
�����B��@-=TF!�QY�}�T�9	�T\���� � �L\��Q�]�w�9M� ��t�b��^�*��7}\x Qb��r�	����G A�w�SP�_��̃�j�j�$� �if��vP��2R�Y�� ��8��JQ��+'lf-�{��Dμ�
Q��jhM4-�/_k��75Cr    IEND�B`� 
BackgroundclWindowNameSave AllPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:54+01:00" xmp:MetadataDate="2022-09-01T11:07:54+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e4c4be3e-672e-ec47-9f06-0e948f0d2018" xmpMM:DocumentID="adobe:docid:photoshop:9e79f5ef-2bf9-484e-bfda-3cafbd57be4b" xmpMM:OriginalDocumentID="xmp.did:d2565718-62cf-2c4d-bd36-daf99c4b79e5"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d2565718-62cf-2c4d-bd36-daf99c4b79e5" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e4c4be3e-672e-ec47-9f06-0e948f0d2018" stEvt:when="2022-09-01T11:07:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���l  �IDATxڭ�MkA�gZ��� ��RiAi��(bAQ?���v�� ^��/
�� 
4&mlm�T-����&"�Ѓ�D�mw�����tg��4����������V	��"B�~!|�l������|�3�϶aJ,7�>�X%�/|_n�E�� �_0�������ε�4�R �O�⭦�Pnҭ�X2h��q��2�M:#R �E�.��H�d�,@��#o�k�Aq���&�LEG�f�3� ��:���H��\�ۛ>w�@`U�n�#�y<@���"Q�b"��9���~������$d�
�_��0-�nBDP�����y���#4\ �?������Ƿ��Y�rw���#� ��?>��&0�v T��1 =����	<�u����T�Y0ҭ\_�2��j�B3ڜ�z�j����%�3\׮uP��t|�_����16�
�^��EV�r�q�����ý��~�@�c�`���h�l��t]��`����`�T�4{�o�3�pݸ������h7�W,��ɲF��)X?b=���4���`VC����äY~�;����ѽ�� Q��`�Kヤɹ�U��t|��v5���!\8{�49_[#�{�8ގ?�f|���.2�,��H�˟����������3���@p�)XL�芃�U3����N%�    IEND�B`�  Left(Top    TPF0TEditorPreferencesDialogEditorPreferencesDialogLeft/Top� HelpType	htKeywordHelpKeywordui_editor_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionEditorPreferencesDialogClientHeight~ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�~ 
TextHeight 	TGroupBoxExternalEditorGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionC   Alternativ extern editor (påverkar bara redigering av fjärrfiler)TabOrder
DesignSize�I  	TCheckBoxExternalEditorTextCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight CaptionH   Tvinga fram textöverföringsläge för filer redigerade i extern editorTabOrder  	TCheckBoxSDIExternalEditorCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionA   E&xtern editor öppnar varje fil i ett separat fönster (process)TabOrder    	TGroupBoxEditorGroup2LeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionEditorTabOrder 
DesignSize��   TRadioButtonEditorInternalButtonLeftTopWidth� HeightCaption&Intern editorTabOrder OnClickControlChange  TRadioButtonEditorExternalButtonLeftTop-Width� HeightCaption&Extern editorTabOrderOnClickControlChange  THistoryComboBoxExternalEditorEditLeftTopDWidth6HeightAutoCompleteAnchorsakLeftakTopakRight TabOrderTextExternalEditorEditOnChangeControlChangeOnExitExternalEditorEditExit  TButtonExternalEditorBrowseButtonLeftVTopCWidthPHeightAnchorsakTopakRight Caption   B&läddra...TabOrderOnClickExternalEditorBrowseButtonClick  TRadioButtonEditorOpenButtonLeftTopaWidth� HeightCaption&Associerad applikationTabOrderOnClickControlChange  TButtonDefaultButtonLeft	TopxWidth� HeightCaption    Använd systemets standardeditorTabOrderOnClickDefaultButtonClick   	TGroupBox	MaskGroupLeftTop� Width�HeightIAnchorsakLeftakTopakRight CaptionAutomatiskt val av editorTabOrder
DesignSize�I  TLabel	MaskLabelLeft	TopWidth� HeightCaption/   Använd den här editorn för &följande filer:FocusControlMaskEdit  THistoryComboBoxMaskEditLeft	Top(Width�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder Text*.*OnExitMaskEditExit   TButtonOkButtonLeft� Top]WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeftTop]WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftgTop]WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  	TCheckBoxRememberCheckLeftTopFWidth�HeightAnchorsakLeftakRightakBottom Caption   &Kom ihåg den här editornTabOrder     TPF0TFileFindDialogFileFindDialogLeftoTop� HelpType	htKeywordHelpKeywordui_findBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionFindXClientHeight�ClientWidth2Color	clBtnFaceConstraints.MinHeight� Constraints.MinWidth�Font.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 	Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                  $$*)&�-+)�1/,�51/�+++                                                                                                                                                                                                                                    (   +)%�.,)�1/-�520�853�<85�+++                                                                                                                                                                                                                            (   +)%�.,)�1/-�520�853�<96�?<8�B>:�                                                                                                                                                                                                                        (   +)%�.,)�1/-�520�853�<96�?<8�B?;�FB=�                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������    (   +)%�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������(   +)%�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LHE�                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������+)%�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LGE�II@                            ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������863�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LGE�HH@                                 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������CA?�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LGE�HH@                                     ������������������������������������������������������������������������������������������������������������������������������������������������������������������������CA@�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LGE�HH@                                         ��������������������������������������������������������������������������������������������������������������������������������������������������������������������CA@�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LGE�HH@                                             ����������������������������������������������������������������������������������������������������������������������������������������������������������������CA@�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LGE�HH@                                                 ������������������������������������������������������������������������������������������������������������������������������������������������������������]\Z�.,)�1/-�520�853�<96�?<8�B?;�FB>�IEB�LGE�HH@                                                     ����������������������������������������������������������������������������������������������������������������������������������������������������������������@><�520�853�<96�?<8�B?;�FB>�IEB�LGE�HH@                                                         ��������������������������������������������������������������������������������������������������������������������������������������������������������������������FC@�<96�?<8�B?;�FB>�IEB�LGE�HH@                                                             ������������������������������������������������������������������������������������������������������������������������������������������������������������������������MJF�B?;�FB>�IEB�LGE�HH@                                                                 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������UQM�IEB�LGE�HH@                                                                     ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`\Y�HH@                                                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            �������������������������������������������������������������������������������������������������������������������������������ܼ�������������������������������������                                                                            ���������������������������������������������������������������������������������������������������������������������������������ٹ���������������������������������                                                                            �������������������������������������������������������������������������������������������������������������������������������������ѿ�����������������������������                                                                            ��������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������г�������������������������                                                                            ���������������������������������������������������������������������������������������������������������������������������������������������¿����������������������                                                                            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������ű���������������������                                                                            �������������������������������������������������������������������������������������������������������������������������������������������������ȭ���������������������                                                                            ��������������������������������������������������������������������������������������������������������������������������������������������������ɫ���������������������                                                                            ���������������������������������������������������������������������������������������������������������������������������������������������������ì���������������������                                                                            ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ���������������������������������������������������������������������������������������������������������������������������������������������������׫�������������������������                                                                            �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ��������������������������������������������������������������������������������������������������������������������������������������������������ׯ�����������������������������                                                                            ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            �������������������������������������������������������������������������������������������������������������������������������������й���������������������������������������������                                                                            �����������������������������������������������������������������������������������������������������������������������������˺�����������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                            �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                            �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                    �����������������������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                        �������������������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                            ���������������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                                �����������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                                    �������������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                                        ���������������������������������������������������������������������������������������������������������������������������������������������������<                                                                                                            �����������������������������������������������������������������������������������������������������������������������������������������������<                                                                                                                �������������������������������������������������������������������������������������������������������������������������������������������<                                                                                                                    ���������������������������������������������������������������������������������������������������������������������������������������<                                                                                                                        �����������������������������������������������������������������������������������������������������������������������������������<                                                                                                                            �������������������������������������������������������������������������������������������������������������������������������<                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �����������������������������     �      �      �      �      �      �      �      ?�      �      ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ��     ?��     ��     ���    ���    ���    ���    ���    ���    ?���    ���    ����   ����   �������������������������������������������(   0   `          �%                                                                                                                                                                                         )'%�-+*�3/.�630U                                                                                                                                                                           )'&�.,*�30.�742�:74�>;8W                                                                                                                                                                   )'&�.,*�30.�742�;85�@=9�DA=�                                                                                                                                                               )'&�.,*�30.�742�;85�@=9�DA=�IEA�                ������������������������������������������������������������������������������������������������������������������������������������       )'&�.,*�30.�742�;85�@=9�DA=�IEA�MHD�                ������������������������������������������������������������������������������������������������������������������������������������   )'&�.,*�30.�742�;85�@=9�DA=�IEA�MHD�+++                ������������������������������������������������������������������������������������������������������������������������������������)'&�.,*�30.�742�<96�@=9�DA=�IEA�MHD�+++                    ��������������������������������������������������������������������������������������������������������������������������������TQO�.,*�30.�742�<96�@=9�DA=�IEA�MHD�+++                        ����������������������������������������������������������������������������������������������������������������������������vus�.,*�30.�742�<96�@=9�DA=�IEA�MHD�+++                            ����������������������������������������������������������������������������������������������������������������������������.,*�30.�742�<96�@=9�DA=�IEA�MHD�+++                                ����������������������������������������������������������������������������������������������������������������������������gdb�742�<96�@=9�DA=�IEA�MHD�+++                                    ��������������������������������������������������������������������������������������������������������������������������������okh�@=9�DA=�IEA�MHD�+++                                        ������������������������������������������������������������������������������������������������������������������������������������wso�IEA�MHD�+++                                            ������������������������������������������������������������������������������������������������������������������������������������:KHC_+++                                                ����������������������������������������������������������������������������������������������������������������������������                                                            �������������������������������������������������������������������������������������������������������������������������                                                            �����������������������������������������������������������������������������������������������������������������������                                                            ���������������������������������������������������������������������������������������������������������ӵ�������������                                                            �������������������������������������������������������������������������������������������������������������ÿ������������
                                                        ��������������������������������������������������������������������������������������������������������������ʳ������������L                                                        ���������������������������������������������������������������������������������������������������������������֧������������{                                                        ����������������������������������������������������������������������������������������������������������������ۤ�������������                                                        �����������������������������������������������������������������������������������������������������������������ܤ�������������                                                        ������������������������������������������������������������������������������������������������������������������ק�������������                                                        �������������������������������������������������������������������������������������������������������������������ī������������`                                                        ����������������������������������������������������������������������������������������������������������������������������������                                                        ������������������������������������������������¿����������������������������������������������������������������Э�������������                                                            ����������������������������������������������������������������������������������������������������������������������������������                                                            �����������������������������������������������������������������������������������������������������������������������������������                                                            ���������������������������������������������������������������������������������������������������������޾�������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            ������������������������������������������������������������������������������������������������������������������������������������                                                            �����������������������������������������������������������������������������������������������������������������������������������<                                                            �������������������������������������������������������������������������������������������������������������������������������<                                                                ���������������������������������������������������������������������������������������������������������������������������<                                                                    �����������������������������������������������������������������������������������������������������������������������<                                                                        �������������������������������������������������������������������������������������������������������������������<                                                                            ���������������������������������������������������������������������������������������������������������������<                                                                                �����������������������������������������������������������������������������������������������������������<                                                                                    �������������������������������������������������������������������������������������������������������<                                                                                        ���������������������������������������������������������������������������������������������������<                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������  �����  �����  �����  �     �      �      �      �      �      �    ?  �      �    �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   ?�  �   �  �   ��  �  ��  �  ��  �  ��  �  ��  ������  ������  ������  ������  (   (   P          @                                                                                                                                                              '!!',)(�0.,�641�+++                                                                                                                                        $$$++)(�1/,�641�;85�A<:�                                                                                                                                    $$$++)(�1/,�641�;85�A=:�EB?�                                                                                                                                $$$++)(�1/,�641�;85�A=:�FB?�JFC�            ������������������������������������������������������������������������������������������������������������    $$$++)(�1/,�641�;85�A=:�FB?�KGB�MFF(            ������������������������������������������������������������������������������������������������������������$$$++)(�1/,�641�;85�A=:�FB?�KGB�MGG+                ������������������������������������������������������������������������������������������������������������+)(�1/,�641�;85�A=:�FB?�KGB�MGG+                    ��������������������������������������������������������������������������������������������������������520�1/,�641�<96�A=:�FB?�KGB�MGG+                        ��������������������������������������������������������������������������������������������������������974�641�<96�A=:�FB?�KGB�MGG+                            ������������������������������������������������������������������������������������������������������������B?<�A=:�FB?�KGB�MGG+                                ����������������������������������������������������������������������������������������������������������������KFC�KGB�MGG+                                    �������������������������������������������������������������������������������������������������������������RMM2MGG+                                        ��������������������������������������������������������������������������������������������������������                                                ������������������������������������������������������������������������������������۹�������������                                                    ���������������������������������������������������������������������������������������Ѽ������������                                                 ������������������������������������������������������������������������������������������������������                                                ��������������������������������������������������������������������������������������������ɴ���������                                                ���������������������������������������������������������������������������������������������ը������������                                            ����������������������������������������������������������������������������������������������٥������������                                             �����������������������������������������������������������������������������������������������ئ������������                                            ������������������������������������������������������������������������������������������������ͩ������������                                            ������������������������������������������������������������������������������������������������������������                                                �����������������������������������������������������������������������������������������������ݯ������������z                                                ��������������������������������������������������������������������������������������������������������������                                                ���������������������������������������������¿������������������������������������������������������������                                                    �������������������������������������������������������������������������������������ۿ���������������������                                                    �����������������������������������������������������������������������������Ǽ�����������������������������                                                    ������������������������������������������������������������������������������������������������������������                                                    ������������������������������������������������������������������������������������������������������������                                                    ������������������������������������������������������������������������������������������������������������                                                    ������������������������������������������������������������������������������������������������������������                                                    �����������������������������������������������������������������������������������������������������������<                                                    �������������������������������������������������������������������������������������������������������<                                                        ���������������������������������������������������������������������������������������������������<                                                            �����������������������������������������������������������������������������������������������<                                                                �������������������������������������������������������������������������������������������<                                                                    ���������������������������������������������������������������������������������������<                                                                        �����������������������������������������������������������������������������������<                                                                                                                                                                                                                                                                                                                                                                                                �����   �����   �����   ����    �      �      �      �      �      �      �   ?   �      �  �   �  �   �  �   �  �   �  �   �   �   �   �   �   �   �   �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  ?�   �  �   �  ��   �����   �����   (       @          �                                                                                                                                  ($$G.,(�51/�;728                                                                                                            %%"K.,)�52/�;85�A>:�        ��������������������������������������������������������������������������������������������    %%"K.,)�52/�;85�B>;�HDA�        ��������������������������������������������������������������������������������������������%%"K.,)�52/�;85�B>;�HDA�MKFj        ����������������������������������������������������������������������������������������{wt�.,)�52/�;85�B>;�HDA�NJEr            ����������������������������������������������������������������������������������������0.+�52/�;85�B>;�HDA�NJEr                ������������������������������������������������������������������������������������HFD�52/�;85�B>;�HDA�NJEr                    ����������������������������������������������������������������������������������������GDA�B>;�HDA�NJEr                        ��������������������������������������������������������������������������������������������LGD�NJEr                            ���������������������������������������������������������������������������������������@@@                                �������������������������������������������������������������������������������������                                    �����������������������������������������������������������������������������������                                    �������������������������������������������������������������������������֬���������                                    ������������������������������������������������������������������������������������                                    �������������������������������������������������������������������������������������                                    �����������������������������������������������������������������������������������������                                ���������������������������������������������������������������������������������������                                    ������������������������������������������������������������������������������Ϭ���������                                    ������������������������������������������������������������������������������������������                                    �������������������������������������������������������������������������������������������                                    ���������������������������������������������������������������������ӽ���������������������                                    ��������������������������������������������������������������������������������������������                                    ��������������������������������������������������������������������������������������������                                    �������������������������������������������������������������������������������������������K                                    ���������������������������������������������������������������������������������������K                                        �����������������������������������������������������������������������������������K                                            �������������������������������������������������������������������������������K                                                ���������������������������������������������������������������������������K                                                    �����������������������������������������������������������������������<                                                        �������������������������������������������������������������������<                                                                                                                                                                                                                                                                                                                    ���������  @�   �  �  �  �  �  �  ?�  �  �  �  �  �  ?�  �  �  �  �  �  �  �  �  �� �� �� �� �� ���������(      0          `	                                                                                                      (&$2/,�;82[                                                                                )'#�2/-�;85�D?<�            ����������������������������������������������������������������_\Y�2/-�;85�D@=�LID�            ����������������������������������������������������������������20-�;85�D@=�MHE�               ������������������������������������������������������������20-�;85�D@=�MHE�                   ������������������������������������������������������������GDA�D@=�MHE�                       ����������������������������������������������������������������plh�                           ���������������������������������������������������������������                            �����������������������������������������������ڰ�������������                            ��������������������������������������������������������������                            ����������������������������������������������������Ǯ���������                            �����������������������������������������������������ū���������                            �����������������������������������������������������������������                            ����������������������������������������������������ڰ�������������                            �������������������������������������������������������������������                            ��������������������������������������������������������������������                            ��������������������������������������������������������������������                            �������������������������������������������������������������������K                            ���������������������������������������������������������������K                                �����������������������������������������������������������K                                    �������������������������������������������������������G                                        ���������������������������������������������������<                                                                                                                                                                                                                                ��� ��� �   �   �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � ? �  � � ��� ��� (      (          �                                                                                      %%"K0.,�;74p        ��������������������������������������������������������{wt�1.,�;85�DA>�        ��������������������������������������������������������30.�;85�EA>�NIGl        ����������������������������������������������������521�;85�EA>�NJEr            ������������������������������������������������SPN�;85�EA>�NJEr                ����������������������������������������������������pmj�zvs�                    ���������������������������������������������������������                    ����������������������������������������Ե�������������                    �������������������������������������������������������                    ��������������������������������������������������������                    ���������������������������������������������������������                    ����������������������������������������������������������                    �����������������������������������������������������������                    ������������������������������������������������������������                    ������������������������������������������������������������                    �����������������������������������������������������������K                    �������������������������������������������������������K                        ���������������������������������������������������K                            �����������������������������������������������<                                                                                                        ��� �   �   �  � 0 � p � p � p � p � p � p � p � p � p � p � p � � �� �� ��� (                 @                                                                      -*'�;85�        ��������������������������������������������GEB�;85�GCA�        ����������������������������������������]\Y�;85�HCA�M@@        ����������������������������������������NKH�VRO�M@@            ��������������������������������Ǽ�������������                ��������������������������������������������                ����������������������������������ب���������                �����������������������������������ڧ���������                ������������������������������������é���������                �����������������¿��������������Ѷ�������������                ������������������������������������������������                ������������������������������������������������                �����������������������������������������������K                �������������������������������������������K                    ���������������������������������������<                                                                                ��  �   �   �  �  �  �  �  �  �  �  �  �  �  �  ��  
KeyPreview	PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnClose	FormCloseOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize2� 
TextHeight 	TGroupBoxFilterGroupLeftTopWidth�HeightzAnchorsakLeftakTopakRight CaptionFilterTabOrder 
DesignSize�z  TLabel	MaskLabelLeft1TopWidth4HeightCaption	&Filmask:FocusControlMaskEdit  TLabelRemoteDirectoryLabelLeft1TopGWidth3HeightCaption   Sö&k i:FocusControlRemoteDirectoryEdit  	TPaintBoxAnimationPaintBoxLeftTopWidth Height   THistoryComboBoxRemoteDirectoryEditLeft1TopYWidthvHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxMaskEditLeft1Top(Width HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextMaskEditOnChangeControlChangeOnExitMaskEditExit  TStaticTextMaskHintTextLeft� Top?Width|Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	  TButton
MaskButtonLeftWTop'WidthPHeightAnchorsakTopakRight Caption	&RedigeraTabOrderOnClickMaskButtonClick   TButtonStartStopButtonLeft�TopWidthlHeightAnchorsakTopakRight Caption&StartXDefault	TabOrderOnClickStartStopButtonClick  TButton
HelpButtonLeft�Top.WidthlHeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelFileViewPanelLeftTop� Width�Height� AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder TIEListViewFileViewLeft Top Width�Height� AlignalClientFullDrag	ReadOnly		RowSelect		PopupMenuFileViewPopupMenuTabOrder 
OnDblClickFileViewDblClickOnEnterControlChangeOnExitControlChange
NortonLikenlOffColumnsCaptionNamnWidthP CaptionKatalogWidthx 	AlignmenttaRightJustifyCaptionStorlekWidthP Caption   ÄndradWidthZ  	ViewStylevsReport	OnCompareFileViewCompareOnContextPopupFileViewContextPopupOnSelectItemFileViewSelectItem   
TStatusBar	StatusBarLeft Top�Width2HeightPanels SimplePanel	  TButtonFocusButtonLeft�Top� WidthlHeightActionFocusActionAnchorsakTopakRight TabOrder  TButton
CopyButtonLeft�TopmWidthlHeightAction
CopyActionAnchorsakRightakBottom TabOrder  TButtonDeleteButtonLeft�Top� WidthlHeightActionDeleteActionAnchorsakTopakRight TabOrder  TButtonDownloadButtonLeft�Top� WidthlHeightActionDownloadActionAnchorsakTopakRight TabOrder  TButton
EditButtonLeft�Top� WidthlHeightAction
EditActionAnchorsakTopakRight Caption	&RedigeraTabOrder  
TPopupMenuFileViewPopupMenuLeft�Top 	TMenuItemFocus1ActionFocusActionDefault	  	TMenuItemN1Caption-  	TMenuItemEdit1Action
EditAction  	TMenuItem	Download1ActionDownloadAction  	TMenuItemDelete1ActionDeleteAction  	TMenuItemN2Caption-  	TMenuItemSelectAllItemActionSelectAllAction  	TMenuItemN3Caption-  	TMenuItemCopyResults1Action
CopyAction   TActionList
ActionListLeft�Top= TActionDeleteActionCaption&Ta bortSecondaryShortCuts.StringsF8 ShortCut.	OnExecuteDeleteActionExecute  TActionFocusActionCaptionF&okus	OnExecuteFocusActionExecute  TActionSelectAllActionCaptionM&arkera alltShortCutA@	OnExecuteSelectAllActionExecute  TAction
CopyActionCaption&Kopiera resultatShortCutC@	OnExecuteCopyActionExecute  TActionDownloadActionCaptionLadda &ner...ShortCutt	OnExecuteDownloadActionExecute  TAction
EditActionCaption	&RedigeraSecondaryShortCuts.StringsCtrl+E ShortCuts	OnExecuteEditActionExecute      TPF0TFileSystemInfoDialogFileSystemInfoDialogLeft@Top� HelpType	htKeywordHelpKeyword	ui_fsinfoBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption#Information om server och protokollClientHeight�ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnShowFormShow
DesignSize�� 
TextHeight TButtonCloseButtonLeftTop�WidthPHeightAnchorsakRightakBottom Cancel	Caption   StängDefault	ModalResultTabOrder  TButton
HelpButtonLeftXTop�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPageControlPageControlLeft Top Width�Height�
ActivePageProtocolSheetAlignalTopAnchorsakLeftakTopakRightakBottom TabOrder OnChangePageControlChange 	TTabSheetProtocolSheetCaption	Protokoll
DesignSize�w  	TGroupBoxHostKeyGroupLeftTop� Width�Height_AnchorsakLeftakRightakBottom Caption$   Nyckelfingeravtryck till värdserverTabOrder
DesignSize�_  TLabelLabel2LeftTopWidth9HeightCaptionAlgoritmFocusControlHostKeyAlgorithmEdit  TLabelLabel3LeftTop-Width1HeightCaptionSHA-256:FocusControlHostKeyFingerprintSHA256Edit  TLabelLabel4LeftTopDWidthHeightCaptionMD5:FocusControlHostKeyFingerprintMD5Edit  TEditHostKeyFingerprintSHA256EditLeftXTop-Width:HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFace	PopupMenuFingerprintPopupMenuReadOnly	TabOrderTextHostKeyFingerprintSHA256EditOnContextPopup(HostKeyFingerprintSHA256EditContextPopup  TEditHostKeyAlgorithmEditLeftXTopWidth:HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextHostKeyAlgorithmEdit  TEditHostKeyFingerprintMD5EditLeftXTopDWidth:HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFace	PopupMenuFingerprintPopupMenuReadOnly	TabOrderTextHostKeyFingerprintMD5EditOnContextPopup(HostKeyFingerprintSHA256EditContextPopup   	TListView
ServerViewLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�  Caption   VärdeWidth�   ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup  	TGroupBoxCertificateGroupLeftTopQWidth�HeightfAnchorsakLeftakRightakBottom CaptionCertifikatets fingeravtryckTabOrder
DesignSize�f  TLabelLabel5LeftTopWidth1HeightCaptionSHA-256:FocusControl CertificateFingerprintSha256Edit  TLabelLabel6LeftTop-Width%HeightCaptionSHA-1:FocusControlCertificateFingerprintSha1Edit  TEdit CertificateFingerprintSha256EditLeftXTopWidth:HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder Text CertificateFingerprintSha256Edit  TButtonCertificateViewButtonLeftTopDWidth� HeightCaption   &Fullständigt certifikatTabOrderOnClickCertificateViewButtonClick  TEditCertificateFingerprintSha1EditLeftXTop-Width:HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFace	PopupMenuFingerprintPopupMenuReadOnly	TabOrderTextCertificateFingerprintSha1EditOnContextPopup(HostKeyFingerprintSHA256EditContextPopup    	TTabSheetCapabilitiesSheetCaption   Möjligheter
ImageIndex
DesignSize�w  	TGroupBox	InfoGroupLeftTop� Width�Height� AnchorsakLeftakRightakBottom Caption   Övrig informationTabOrder
DesignSize��   TMemoInfoMemoLeft	TopWidth�HeightfTabStopAnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneColor	clBtnFaceLines.StringsInfoMemo 
ScrollBarsssBothTabOrder WordWrap   	TListViewProtocolViewLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�  Caption   VärdeWidth�   ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupControlContextPopup   	TTabSheetSpaceAvailableSheetCaption   Tillgängligt utrymme
ImageIndex
DesignSize�w  TLabelLabel1LeftTopWidthHeightCaption
   &Sökväg:FocusControlSpaceAvailablePathEdit  	TListViewSpaceAvailableViewLeftTop"Width�Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionArtikelWidth�  Caption   VärdeWidth�   ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupControlContextPopupOnCustomDrawItem SpaceAvailableViewCustomDrawItem  TEditSpaceAvailablePathEditLeft8TopWidth� HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChangeOnEnterSpaceAvailablePathEditEnterOnExitSpaceAvailablePathEditExit  TButtonSpaceAvailableButtonLeft4TopWidthmHeightAnchorsakTopakRight CaptionKon&trolleraTabOrderOnClickSpaceAvailableButtonClick    TButtonClipboardButtonLeftTop�Width� HeightAnchorsakLeftakBottom Caption&Kopiera till urklippTabOrderOnClickClipboardButtonClick  
TPopupMenuListViewMenuLeft� Topb 	TMenuItemCopyCaptionK&opieraOnClick	CopyClick   
TPopupMenuFingerprintPopupMenuLeft� Topb 	TMenuItemCopy1ActionEditCopyAction  	TMenuItem ActionEditSelectAllAction   TActionListFingerprintActionListLeftHTopb 	TEditCopyEditCopyActionCategoryEditCaptionK&opieraShortCutC@	OnExecuteEditCopyActionExecuteOnUpdateEditCopyActionUpdate  TEditSelectAllEditSelectAllActionCategoryEditCaption&Markera alltShortCutA@    TPF0TFullSynchronizeDialogFullSynchronizeDialogLeftmTop� HelpType	htKeywordHelpKeywordui_synchronizeBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynkroniseraClientHeight�ClientWidthColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize� 
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidthHeightxAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSizex  TLabelLocalDirectoryLabelLeft1TopWidthQHeightCaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft1TopEWidth^HeightCaption   F&järrka&talog:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	  THistoryComboBoxRemoteDirectoryEditLeft1TopWWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeft1Top(WidthvHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeft�Top'WidthPHeightAnchorsakTopakRight Caption   Bl&äddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButtonOkButtonLeftTop�Width^HeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrderOnClickOkButtonClickOnDropDownClickOkButtonDropDownClick  TButtonCancelButtonLefthTop�WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder	  	TGroupBoxOptionsGroupLeftTop� Width� HeightyCaption   Alternativ för synkroniseringTabOrder
DesignSize� y  	TCheckBoxSynchronizeDeleteCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeftTop[Width� HeightAnchorsakLeftakTopakRight CaptionBara &valda filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeftTopDWidth� HeightAnchorsakLeftakTopakRight Caption&Endast existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizePreviewChangesCheckLeftTop-Width� HeightAnchorsakLeftakTopakRight Caption   Fö&rhandsvisa ändringarTabOrderOnClickControlChange   TButtonTransferSettingsButtonLeftTop�Width� HeightAnchorsakLeftakBottom Caption   Överf&öringsinställningar...TabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxDirectionGroupLeftTop� WidthHeight1AnchorsakLeftakTopakRight Caption   Riktning/målkatalogTabOrder TRadioButtonSynchronizeBothButtonLeftTopWidth� HeightCaption   &BådaChecked	TabOrder TabStop	OnClickControlChange  TRadioButtonSynchronizeRemoteButtonLeft� TopWidth� HeightCaption   &FjärrTabOrderOnClickControlChange  TRadioButtonSynchronizeLocalButtonLeftSTopWidth� HeightCaption&LokalTabOrderOnClickControlChange   	TGroupBoxCompareCriterionsGroupLeftTop� Width� HeightyAnchorsakLeftakTopakRight Caption   JämförelsekriterierTabOrder
DesignSize� y  	TCheckBoxSynchronizeByTimeCheckLeftTopWidth� HeightAnchorsakLeftakTopakRight Caption   Ä&ndringstidTabOrder OnClickControlChange  	TCheckBoxSynchronizeBySizeCheckLeftTop-Width� HeightAnchorsakLeftakTopakRight CaptionF&ilstorlekTabOrderOnClickControlChange  	TCheckBoxSynchronizeCaseSensitiveCheckLeftTop[Width� HeightAnchorsakLeftakTopakRight Caption   Sk&riftlägeskänsligTabOrderOnClickControlChange  	TCheckBoxSynchronizeByChecksumCheckLeftTopDWidth� HeightAnchorsakLeftakTopakRight CaptionKo&ntrollsummaTabOrderOnClickControlChange   	TCheckBoxSaveSettingsCheckLeftTopsWidth�HeightAnchorsakLeftakTopakRight Caption   Använd &samma val nästa gångTabOrder  	TGroupBoxCopyParamGroupLeftTop�WidthHeight;AnchorsakLeftakTopakRight Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize;  TLabelCopyParamLabelLeft	TopWidth�Height#AnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamGroupClick   TButton
HelpButtonLeft�Top�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrder
OnClickHelpButtonClick  	TGroupBox	ModeGroupLeftTop� WidthHeight1AnchorsakLeftakTopakRight Caption   LägeTabOrder TRadioButtonSynchronizeFilesButtonLeftTopWidth� HeightCaptionSynkronisera &filerTabOrder OnClickControlChange  TRadioButtonMirrorFilesButtonLeft� TopWidth� HeightCaptionS&pegelfilerTabOrderOnClickControlChange  TRadioButtonSynchronizeTimestampsButtonLeftSTopWidth� HeightCaption   Synkronisera tidss&tämplarTabOrderOnClickControlChange   
TPopupMenuOkMenuLeft�Top� 	TMenuItemStart1Caption&StartDefault	OnClickStart1Click  	TMenuItemStartInNewWindowItemCaption   Starta i &nytt fönsterOnClickStartInNewWindowItemClick       TPF0TGenerateUrlDialogGenerateUrlDialogLeftqTopHelpType	htKeywordHelpKeywordui_generateurlBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionGenerate URL XClientHeight}ClientWidthColor	clBtnFaceConstraints.MinHeight,Constraints.MinWidth�Font.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnShowFormShow
DesignSize} 
TextHeight TPageControlOptionsPageControlLeft Top WidthHeighth
ActivePageUrlSheetAnchorsakLeftakTopakRight TabOrder OnChangeControlChange 	TTabSheetUrlSheetCaptionURL 	TCheckBoxUserNameCheckTagLeftTopWidth� HeightCaption   &AnvändarnamnTabOrder OnClickControlChange  	TCheckBoxHostKeyCheckTagLeft� TopWidth� HeightCaption   SSH &värdnyckelTabOrderOnClickControlChange  	TCheckBoxWinSCPSpecificCheckTagLeft� TopWidth� HeightCaptionWinSCP-specifikTabOrderOnClickControlChange  	TCheckBoxSaveExtensionCheckTag Left� Top3Width� HeightCaption   &Spara sessionsinställningarTabOrderOnClickControlChange  	TCheckBoxRemoteDirectoryCheckTagLeftTop3Width� HeightCaptionInitial &katalogTabOrderOnClickControlChange  	TCheckBoxPasswordCheckTagLeftTopWidth� HeightHelpType	htKeywordCaption
   &LösenordTabOrderOnClickControlChange  	TCheckBoxRawSettingsCheckTag@LeftATopWidth� HeightCaption   &Avancerade inställningarTabOrderOnClickControlChange   	TTabSheetScriptSheetCaptionSkript
ImageIndex
DesignSizeJ  TLabelLabel2LeftTopWidth)HeightCaption&Format:FocusControlScriptFormatCombo  TLabelScriptDescriptionLabelLeftTop WidthHeight*AnchorsakLeftakTopakRightakBottom AutoSizeCaptionScriptDescriptionLabelShowAccelCharWordWrap	  	TComboBoxScriptFormatComboLeftjTopWidth� HeightStylecsDropDownListTabOrder OnChangeControlChangeItems.Strings	SkriptfilBatchfilKommandoradPowerShell-skript    	TTabSheetAssemblySheetCaption.NET assemblerkod
ImageIndex
DesignSizeJ  TLabelLabel1LeftTopWidth7HeightCaption   &SpråkFocusControlAssemblyLanguageCombo  TLabelAssemblyDescriptionLabelLeftTop WidthHeight*AnchorsakLeftakTopakRightakBottom AutoSizeCaptionAssemblyDescriptionLabelShowAccelCharWordWrap	  	TComboBoxAssemblyLanguageComboLeftjTopWidth� HeightStylecsDropDownListTabOrder OnChangeControlChangeItems.StringsC#VB.NET
PowerShell     	TGroupBoxResultGroupLeftTopnWidthHeight� AnchorsakLeftakTopakRightakBottom CaptionResultXTabOrder
DesignSize�   TMemo
ResultMemoLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneTabOrder    TButton	CancelBtnLeftmTop\WidthPHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  TButton
HelpButtonLeft�Top\WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClipboardButtonLeftTop\Width� HeightAnchorsakLeftakBottom Caption&Kopiera till urklippTabOrderOnClickClipboardButtonClick   TPF0TImportSessionsDialogImportSessionsDialogLeftjTop� HelpType	htKeywordHelpKeyword	ui_importBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionImport sitesXClientHeight3ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnShowFormShow
DesignSize�3 
TextHeight TLabelLabelLeftTopWidthDHeightCaption   &Importera från:FocusControlSourceComboBox  TButtonOKButtonLeft� TopWidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� TopWidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  	TListViewSessionListView2LeftTop'Width�Height� AnchorsakLeftakTopakRightakBottom 
Checkboxes	ColumnsWidth�   ColumnClickDoubleBuffered	HideSelectionReadOnly	ParentDoubleBufferedParentShowHintShowColumnHeadersShowHint	TabOrder	ViewStylevsReport	OnInfoTipSessionListView2InfoTipOnKeyUpSessionListView2KeyUpOnMouseDownSessionListView2MouseDown  TButtonCheckAllButtonLeftTopWidth}HeightAnchorsakLeftakBottom CaptionMarkera/avmarkera &allaTabOrderOnClickCheckAllButtonClick  TButton
HelpButtonLeftJTopWidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  	TComboBoxSourceComboBoxLefttTop	Width� HeightStylecsDropDownListTabOrder OnSelectSourceComboBoxSelectItems.StringsPuTTYKiTTY	FileZillaOpenSSHINI fileknown_hosts   TPanel
ErrorPanelLeft0Top\WidthAHeight}
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder TLabel
ErrorLabelLeft Top WidthAHeight}AlignalClient	AlignmenttaCenterCaption
ErrorLabelShowAccelCharLayouttlCenterWordWrap	   TButtonPasteButtonLeft� TopWidthKHeightCaptionKl&istra inTabOrderOnClickPasteButtonClick  TButtonBrowseButtonLeft� TopWidthPHeightCaption   Blädd&ra...TabOrderOnClickBrowseButtonClick    TPF0TLicenseDialogLicenseDialogLeft�Top� ActiveControlCloseButtonBorderIconsbiSystemMenu BorderStylebsDialogCaption   AnvändarlicensClientHeightcClientWidth/Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenter
DesignSize/c 
TextHeight TButtonCloseButtonLeft�TopBWidthPHeightAnchorsakRightakBottom Cancel	Caption   StängDefault	ModalResultTabOrder   TMemoLicenseMemoLeftTopWidthHeight4AnchorsakLeftakTopakRightakBottom Color	clBtnFaceReadOnly	
ScrollBars
ssVerticalTabOrderWantReturns   TPF0TLocationProfilesDialogLocationProfilesDialogLeftWTop� HelpType	htKeywordHelpKeywordui_locationprofileBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionPlatsprofilerClientHeight�ClientWidthYColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnShowFormShow
DesignSizeY� 
TextHeight TLabelLocalDirectoryLabelLeft.TopWidthQHeightCaptionL&okal katalog:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft.Top7Width^HeightCaption   F&järrkatalog:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	  TButtonOKBtnLeftUTop�WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft�Top�WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTopfWidthIHeight3
ActivePageSessionProfilesSheetAnchorsakLeftakTopakRightakBottom TabOrder 	TTabSheetSessionProfilesSheetTagCaptionSessionsplatsprofiler
DesignSizeA  	TTreeViewSessionProfilesViewTagLeftTopWidth�Height
AnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionIndentParentDoubleBufferedTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDragItems.NodeData
                ��������           1 "           ��������            1 1             ��������            2             ��������            3            ��������           4 "           ��������            4 1             ��������            5   TButtonAddSessionBookmarkButtonTagLeft�TopWidth\HeightAnchorsakTopakRight Caption   &Lägg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeft�Top$Width\HeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeft�Top� Width\HeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�Left�Top� Width\HeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonRenameSessionBookmarkButtonTagLeft�TopCWidth\HeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSessionBookmarkMoveToButtonTagLeft�TopbWidth\HeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick   	TTabSheetSharedProfilesSheetTagCaptionDelade platsprofiler
ImageIndex
DesignSizeA  	TTreeViewSharedProfilesViewTagLeftTopWidth�Height
AnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionImagesBookmarkImageListIndentParentDoubleBufferedTabOrder OnChangeProfilesViewChangeOnCollapsedProfilesViewCollapsed
OnDblClickProfilesViewDblClick
OnDragDropProfilesViewDragDrop
OnDragOverProfilesViewDragOverOnEditedProfilesViewEdited	OnEditingProfilesViewEditing	OnEndDragProfilesViewEndDrag
OnExpandedProfilesViewExpandedOnGetImageIndexProfilesViewGetImageIndexOnGetSelectedIndexProfilesViewGetSelectedIndex	OnKeyDownProfilesViewKeyDownOnStartDragProfilesViewStartDragItems.NodeData
                ��������           1 "           ��������            1 1             ��������            2             ��������            3            ��������           4 "           ��������            4 1             ��������            5   TButtonAddSharedBookmarkButtonTagLeft�TopWidth\HeightAnchorsakTopakRight Caption   &Lägg till...TabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeft�Top$Width\HeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonRenameSharedBookmarkButtonTagLeft�TopCWidth\HeightAnchorsakTopakRight Caption	B&yt namnTabOrderOnClickRenameBookmarkButtonClick  TButtonSharedBookmarkMoveToButtonTagLeft�TopbWidth\HeightAnchorsakTopakRight Caption&Flytta till...TabOrderOnClickBookmarkMoveToButtonClick  TButtonUpSharedBookmarkButtonTag�Left�Top� Width\HeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeft�Top� Width\HeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeft�Top� Width\HeightAnchorsakTopakRight Caption   &Genväg...TabOrderOnClickShortCutBookmarkButtonClick    THistoryComboBoxLocalDirectoryEditLeft.TopWidth�HeightAnchorsakLeftakTopakRight DropDownCountTabOrder TextLocalDirectoryEditOnChangeDirectoryEditChangeSaveOn   THistoryComboBoxRemoteDirectoryEditLeft.TopIWidth#HeightAnchorsakLeftakTopakRight DropDownCount	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeDirectoryEditChangeSaveOn   TButtonLocalDirectoryBrowseButtonLeftTopWidthPHeightAnchorsakTopakRight Caption   Blädd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop�WidthaHeightAnchorsakLeftakBottom Caption   &Bokmärken...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeftTop�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPngImageListBookmarkImageList	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
5  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:01+01:00" xmp:MetadataDate="2022-09-01T11:02:01+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:116e451d-46f3-db48-9bee-957f8c8366a8" xmpMM:DocumentID="adobe:docid:photoshop:f6cec39b-2e3e-5d47-a939-d81c075fba5d" xmpMM:OriginalDocumentID="xmp.did:43f7417e-d11e-e145-99b0-8e5410fb7efd"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:43f7417e-d11e-e145-99b0-8e5410fb7efd" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:116e451d-46f3-db48-9bee-957f8c8366a8" stEvt:when="2022-09-01T11:02:01+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>Vu��  IDATx�c���?%���N!Y&� �?_ZO�:�����'-���&b�}����g�@l�Ō�wK�2�P���0���YΫD�pF&�%@y�ĳ��<� 7��n)�~��?�����d�b,��(���e�{5��{`>o�n 3�8×����CH���f����W.��<`^l3���%
t�?�$3��6����.C��R�j�202�30(V2��s����X8��`��g`����U�n��e�!�������Ā�k��K�D001���4�X�~�{� �41�����]�WJ��5L����?�j@� X3H��$�#Q��_��C3�bЫ�.O��A$�΃{a�T�Y�a�hy����W�n� ��g����(�j�CTR�� "�����Ci�0��4#��_��3$@��m~o�VH]gd��	������v���r�?������� kb`�%�4���Dʭ}��~"*���jDV�$q �� ��8    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:08+01:00" xmp:MetadataDate="2022-09-01T11:06:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5f0285a2-1a20-234b-9a43-8da79e79cb07" xmpMM:DocumentID="adobe:docid:photoshop:9a4cfe93-5052-9246-bf53-fd91397c86e1" xmpMM:OriginalDocumentID="xmp.did:ed00465a-0d10-4b4e-a04b-d555174bc285"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ed00465a-0d10-4b4e-a04b-d555174bc285" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5f0285a2-1a20-234b-9a43-8da79e79cb07" stEvt:when="2022-09-01T11:06:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Z��  �IDATxڭS9KQ���l�V�PW#*Z��I�Bk� Z��o�j����^�Q�� o���&;Ƹ� t�ͼ���73���3��V���T c�q)p5�;�U%�46�=���vI'��C���T�����?URq�Ͽ���I[Q�8G����X�*A�N8��Y���۲�B�R��W��`����+`j@\KZ�,$y���~�:�����3� `;p����(���iTF]k��JГ���8��ȼa������S	vDdj�^x�����$l��iSϪ�IS�t��{�|�����֮�<լqr��	)p��7;K�Q�؞�Z�8������j�v����Cy�l�ai"==L��Q[����)����Q^�~�@�F����_�� &M?�ZP    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:06+01:00" xmp:MetadataDate="2022-09-01T11:02:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:72f8666d-2ee5-344b-aa1d-a1c6ea8cd32b" xmpMM:DocumentID="adobe:docid:photoshop:cba89235-7918-cb4d-9b5c-ca3e0435cf2a" xmpMM:OriginalDocumentID="xmp.did:7bb19fbd-fb7b-5f47-87b8-73ea5303e6e4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7bb19fbd-fb7b-5f47-87b8-73ea5303e6e4" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:72f8666d-2ee5-344b-aa1d-a1c6ea8cd32b" stEvt:when="2022-09-01T11:02:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��t�  mIDATx�c���?%���N!Y&� �?_ZO�:�����F�Ō�wK�2�Pe���=�!ʀ_����P���?�=�r��;� �1~ކ� fNqf.i �� ���������\N�y���f���K�j�$3��6���oH�����������X�6��ݮ����a`��*�����{������4�����fje�91��Z���:L��!
�h���r��4��]�WJ��5L���M3�fuy�d�~$A(.z���)� � �6��P��"�g�8T3���5�h���NP��j����4���Q5��6�7Ԁ+��32��d~$:20ܒ{
�+��fg }6�e>M    IEND�B`�  Left`Top�   TPngImageListBookmarkImageList120HeightWidth	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:02+01:00" xmp:MetadataDate="2022-09-01T11:02:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:72b73e50-dff1-f34d-a0f8-2bfe5d980132" xmpMM:DocumentID="adobe:docid:photoshop:228dafde-a445-a84f-9b85-b1bd22bd94ae" xmpMM:OriginalDocumentID="xmp.did:cfc306e0-350b-804b-952b-f1e2637223ac"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cfc306e0-350b-804b-952b-f1e2637223ac" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:72b73e50-dff1-f34d-a0f8-2bfe5d980132" stEvt:when="2022-09-01T11:02:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�^��  �IDATx���?lQ��;��ǣ�Ҵi��'�i����bL��8�jb�i\��X�L\��1qҡqk��&�iR
FZ*mE�-(���=���q�:��.�w���>�~�w@(�����`)��r��'LR�ǽ�/��0$y�[�=�)���t?Y^l������7v���Q<�8�6!_��}E	o�I{�o����ySz�8�٫���SE�')�|�L������_�����]���ݳvB�*)H�l��Z���1��z�P�W����� x���s�OF4�6�#���,�����/ݧT��lq*oU�:he(eP��Q��� �A���Dv�N�i3�>�7r!J��J�8˱
�t)�!j,;�@�\y�ޣ7� �@y,.�10�l���28�l ����kqa��n�8��&xj� <|����-Ƴ��V�C��yVsC�s�BK��`9�C��4�1
�k`�>�ծ=m1��H�	�88��x�����rb��:��s��84�a(��т.e4�v{�Y}��*=����$�(�.�~�C魄�~��)��Xw�m���	B([���I�އ��'�I���I]t��W怤���DH�Nm)��D���Ԇ�w:伲����Ƽ���'un��A��    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:09+01:00" xmp:MetadataDate="2022-09-01T11:06:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c9283f14-3d59-ec42-94c8-a53f7ac56617" xmpMM:DocumentID="adobe:docid:photoshop:39bb9190-aaa7-5f45-8ad3-4816d448e4c3" xmpMM:OriginalDocumentID="xmp.did:8f445be8-9da7-1a46-99ef-30686812fd01"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8f445be8-9da7-1a46-99ef-30686812fd01" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c9283f14-3d59-ec42-94c8-a53f7ac56617" stEvt:when="2022-09-01T11:06:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��Q5  �IDATx��MOA�����R���z��F�Ҙ� B?��iL<y ��K4�WCԛH0��Xhm�����<l���mnN��ϼ<��?��#"\fc�)��ap��	P�=�3�//|k+�&	��M���Z�Rb���7��b
��Ѱ�j���"zo'��r��=+�I�A>(S�B�9����:�KV./��F]�:��j�Ջ�� ֑c���A��S%��q��_��?�u`I�
�igAE.�'�A��r��y	<~�oʼ���[��������f�eF%���UY7v�8�d����v�A�L��ԇ�F$��&F'4��#ݸ�|L��-��l`�|�N~}*��5�
�~�)�E����_0ތ��_��ΒV��
���9�~n��U��q<2�sOWG�G��xz�-��g����g���I�.��]������~ReI���{���a�1�D�Ѷ���V���������˫�ҵ�v=���ul�L.��l�pP�q�r{    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:07+01:00" xmp:MetadataDate="2022-09-01T11:02:07+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:97d12c2e-ed65-a447-958b-fe256ac98664" xmpMM:DocumentID="adobe:docid:photoshop:469e9482-7664-3f42-92cf-ba17ffa1700a" xmpMM:OriginalDocumentID="xmp.did:62777e29-adc1-d44f-acc9-9c4ebedb8b10"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:62777e29-adc1-d44f-acc9-9c4ebedb8b10" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:97d12c2e-ed65-a447-958b-fe256ac98664" stEvt:when="2022-09-01T11:02:07+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>6�L  �IDATx�c���?5��0��.aY&d	����|u����!C�6���@!!L�S�ܞ�l��=��������Ny�wٝ_�#�@&qFi ����Q��_~e��̃b����Y9� ���Ҍ,���<r�C�����P�����A��������������] j;�п��g`������@�?�f�ߟ63!��T��S�/�����V��/B!>�pV�[�>Z%�_�8��M.>̥�N�h����k���.O�����ho���2��x�	������:�a�������*v�<��Q�����$~�j8��~c�&���� m*��L������e��0�0���|�R�:#��O@�GB%: �tK6�i��� ����0    IEND�B`�  Left`Top�   TPngImageListBookmarkImageList144HeightWidth	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
R	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:02+01:00" xmp:MetadataDate="2022-09-01T11:02:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:50e6f73d-e067-db41-8b94-ebe9b006364f" xmpMM:DocumentID="adobe:docid:photoshop:7857c06d-4ace-c940-939d-89bf5ce1453a" xmpMM:OriginalDocumentID="xmp.did:e67e81f8-8451-bd4d-9f94-8e2f5f22b037"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e67e81f8-8451-bd4d-9f94-8e2f5f22b037" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:50e6f73d-e067-db41-8b94-ebe9b006364f" stEvt:when="2022-09-01T11:02:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�F  /IDATx�ݕKOQ��g��� 	Bb��@1��Fa!����ct�DE�Q�_A���.�jtA�4�&��ąiA�X�mi��v:�;���a@\��$��=����s�� �1�KC�`�.b���w���"�$���cB��`n\q�+���D�,�S�TI+ �g������/[;S���Po�#D�b�~٣��R������3J��{�&5�PK���	�T�$�}�8�z� �pVH�X ��I���f������#lی��y7v4[���'�������ww��F*
��� �/���� �5d�2����R� K9��F���	P ��w)ْ�R�ˀi�Ѐ%o3.�l#_���I������)	�,D<����E��Ƕ�р�g\�xK�/D��2&)�@ +C�������$�sM� _/��d��ڗ�ϓ
�j f��myq������B%��$������*"	�!��9��K�Z%(�i�H ���|~������h�U>���` [+��Ò��8��ڢת�?D �i@��Q.Y���OS��*!�L � ��L��xA\Ӫ�O���7D��:���`O���POQ*��Ef'��������l%Y�q�=��/�@x������j�d,�ٲ��� b���g����*���W40<�t+g`m3��WKO�q`���>��B��Ukb	���@N6D~˒G�;AGM���X��A��� ![��������HG?�)x����H�`�G�U@����0Z�&�$�	���e�y}��7C\�3#    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:10+01:00" xmp:MetadataDate="2022-09-01T11:06:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:fd6e66cb-f739-d84c-95b7-eef321ba62df" xmpMM:DocumentID="adobe:docid:photoshop:7f4f77c0-967a-ec4e-b48e-be0adc9f4ead" xmpMM:OriginalDocumentID="xmp.did:0f2d0182-2614-614c-8d72-1d030f1ed156"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:0f2d0182-2614-614c-8d72-1d030f1ed156" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:fd6e66cb-f739-d84c-95b7-eef321ba62df" stEvt:when="2022-09-01T11:06:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�,�>  �IDATx���kQƿ�Wk$��Q�LJD�Y1mƅP""�&�U� 1�\������?ЅQ[�
"�R7)��G ڔ6jZL��dr���i2�W�Bw��93�~���9�aD��<��%@�u`�����(s���wK��I�m��@�Y�i�\aU����s0/Xʓ1��_�<AV��[6�ȠX�w��#8	�wo�P�ˬ
�^	�N����s([��Ȃ�u�y�S�F�@z��'���/5@�u�k����ϼ!.b$�U�� j��MPz� Dfu��1��=XS�O��B���u7�JT��) ư�����۰�����X��Q��_�G��Hb���'��M�r	�b2�z����FL;�|����y %އC�[r� vwc�YU�q���T@�@+~x����f�T�䦱sFҔk��
��
R����.����Z�������X&��}[�H4��M)��n�& �����/��:I��Ñ�K�J�7��W�g��*2Oƈ�����x��J�i@��{�X�F���0�Cax}�źo�P�W/��[~V|}&�{ CN(����hvpCee��>�&!��G�}��r��?�R�W�v��%L�z'����ʝ0    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
/  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:08+01:00" xmp:MetadataDate="2022-09-01T11:02:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8dcc1edf-ea10-fe40-999a-4a132ce4705f" xmpMM:DocumentID="adobe:docid:photoshop:70aad4b4-afab-094d-89a9-98dd4e7b2aa4" xmpMM:OriginalDocumentID="xmp.did:cf0fee2a-b160-df41-88f2-e5159d137eb0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cf0fee2a-b160-df41-88f2-e5159d137eb0" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8dcc1edf-ea10-fe40-999a-4a132ce4705f" stEvt:when="2022-09-01T11:02:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>D��  IDATx�ݔOKA��Yvmڨ�L{i)�=�E��"RJ�ԃ�$Ń�A���~<��` '��{(�#=c�l���f�;���!�]ޝy~����D�~r? ��D]Z�=�
�)m���T�7m�|<�n��|�V?�Z�3�y�ω�w��,�-�B��E���.� �Z�!@xܴ��i?w.��l\�WŴ �����EPcl5\A^]6�y�G@��	�%@QC���d�hOA(��bl���`�Nu��k
�RY8׹%J.C8:�q�Z֫��%G )'�����.��	|��c��LF۝_�.����)�o�B�����։J��� �8|˜s��ۍ��$�~t�{����ڴ[��!�D����!��Q���3��uφ��9| /�p&F �	Qy�0�����r]8��x������h/�oGu�c�S��������Q2nh��a;5����V�4�r��oK���D�DQ���h����(��~����܏���;    IEND�B`�  Left`Top  TPngImageListBookmarkImageList192Height Width 	PngImages
BackgroundclWindowNameBookmarkPngImage.Data
�	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:03+01:00" xmp:MetadataDate="2022-09-01T11:02:03+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:865b0991-cb42-1545-918e-c8a0731a8792" xmpMM:DocumentID="adobe:docid:photoshop:e9c8dbf3-eda8-2b4f-b843-9c032cf11826" xmpMM:OriginalDocumentID="xmp.did:8d6a3bbd-9685-cc48-a2db-78cdceb0f445"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8d6a3bbd-9685-cc48-a2db-78cdceb0f445" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:865b0991-cb42-1545-918e-c8a0731a8792" stEvt:when="2022-09-01T11:02:03+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��}  qIDATx��]HQ�ϝu\�u3�u�E�@--�Q!"J��~�@!�]K����z�zz��1�������o��C�5����������W����9s�=�=��Ac��m l �7 ��ԁQDE��0ƽ��ٞ�8�o8*�9�. ���]���^TCQ��P�L��?���˫�C��r�Eba%��e���d���W܏Z�A���'� i,�KB
yV++�a����sw��2�@g9�3�e��kDݼ�WE_������8���VM J����Z��V�=8��o�[��9f�h�m����z��T
T�2��p#֛l�a��L98��O�KS\0��,��c�� K��@w�=`�A!.���-��#;�81��gy�9 �n�D�S}&Lݷr �	1�܃Es��yIȵ[%6��чG5 �;%x#a�ZP>�
�9�\����k �s(v�e!�ͱ����\��x�b�tݤ����!�r(/����m�(�t����sR�]����aF� ��,I�"�D׻4 ��D;d�'�%�x�*)�L��0/��}Vz�age��|$G�n�Bq�6��3�|�:B)z�/* ���hhX+O*�ΉP�R�u��8���'PqBq�,�J���#M!��y\�_ �����F0_H_#���C���bPn�$�a� eMI���Rt13D��Nc� �����/�d�1���.&t�B�CAWF� ށ
l0�!3�[4�����\N/�F�T���"��-�&�s?ךnnQM��kˡ#��X>��? eS�Z�!�~��a��6%EzB��l�f�=!Bh.�c�ɸb٪�O�"�_�R�u4��dЯ��v��;j�������p���ҍ� � �����:    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
e	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:10+01:00" xmp:MetadataDate="2022-09-01T11:06:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6123b322-6c8d-8647-8f82-86944185aaea" xmpMM:DocumentID="adobe:docid:photoshop:49750230-1405-654a-b5b3-f7b1a60aa2fc" xmpMM:OriginalDocumentID="xmp.did:5a3be35d-af8f-444f-b58f-3c89f571b4af"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5a3be35d-af8f-444f-b58f-3c89f571b4af" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6123b322-6c8d-8647-8f82-86944185aaea" stEvt:when="2022-09-01T11:06:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>x���  BIDATx��KLQ���k�-��}h��(�� A��F��L�ׂ�;��r�J�#nLt�EY�R�1�B�P���vǙi;L;3ehH�L��̝����AD(d#��� ���ҏ@�� �pW�����E f��j�g��Ku����s�!�����?f
 �(�H'�O�D�� ßnX�.�@�Q=b�����2��5j�4VZr(HT�R�+���PT�@Uª[<<��"@�2�b��h��(�ʛ�������a�@�����ъkX ��ER�.,��0-�Ė@$��]���Vh� �/dZ).�B�;ll�_,� ���&?������jPE@�'�F\��~s��"���$ �oG_�Z����%�+M�Y�(D8FʆW)�g1QG��	� �gI�����F��ڗ���@�JQ%�u�xr<�Č��Cz
~?M�F�P����W�H��^�U��!S�{���I҄3&��~�le��ʒ�J6��q�,�O����n�?6@sϥ�"�N�5��d	3��iOq���0�ȍ1��հ��X����!��?e�{2v��C7�狡һ�;�5ͣQsz��" 1d���� ��qra���-E:�Nk���i�E ��������N��R��yV�D�4��-8��@�^[5x|���
L���N�6�2�Eg�XW�)/�k��-�;�����[U��q�C�{�JI2<��98N�( >߭A��6(-�����l�Z/,���?-��( ��o��m��|����9Dr�s��7a![��FH��ɔ��    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
l  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:08+01:00" xmp:MetadataDate="2022-09-01T11:02:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e7bbcac2-09c2-9741-bba9-a721dd2243cb" xmpMM:DocumentID="adobe:docid:photoshop:d839a3d1-87ad-2f49-98b3-f353c535cb1b" xmpMM:OriginalDocumentID="xmp.did:733049d7-dcc9-644f-864b-ee70f7c2ee15"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:733049d7-dcc9-644f-864b-ee70f7c2ee15" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e7bbcac2-09c2-9741-bba9-a721dd2243cb" stEvt:when="2022-09-01T11:02:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  IIDATx�c���?�@�Q�:`P8��^�	��r�302aU������v�絔X�ͳ`��#���(0�:b-��{�4Q� �w?����~�b@@.`d���?#�TV�g9��[��Y:�����T�3��p��I{:#V��,��LL��b��?��3ÿ?@s���06���ȁ���W��Io	v����W��G{Z�������5�r�e��B�cd���l{	����/k^�Є�d������� |����h����H���b�r�`�Y��Q����8�,��a���(V�{x`��#(��o��EOt�e�:?�� �t�f9������<0J��j�9
��X]��q�a�
W�b�A���bQ�yS����w�~$�Fl���G�!���ð #(Iu���Q��_<Y��F���:�Dd+\�B+���xh�,ˉsv�	;@Ӄ���?�:< � ��v=q�?�T��<�ܢ�W���_��#�R���>8�@zP&���19 �&���raO�:` ��;  �� �h��s    IEND�B`�  Left`Top@   TPF0TLoginDialogLoginDialogLeft_Top� HelpType	htKeywordHelpKeywordui_loginBorderIconsbiSystemMenu
biMinimizebiHelp Caption
InloggningClientHeight�ClientWidthiColor	clBtnFaceConstraints.MinHeight�Constraints.MinWidth�Font.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 
KeyPreview	PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnCloseQueryFormCloseQueryOnShowFormShow
TextHeight TPanel	MainPanelLeft�Top Width�Height�AlignalRight
BevelOuterbvNoneTabOrder  TPanelContentsPanelLeft Top Width�HeightaAlignalClient
BevelOuterbvNoneTabOrder Visible
DesignSize�a  	TGroupBoxContentsGroupBoxLeftTopWidth�HeightVAnchorsakLeftakTopakBottom CaptionContentsGroupBoxTabOrder 
DesignSize�V  TLabelContentsLabelLeftTopWidth#HeightCaptionNamn:ShowAccelChar  TEditContentsNameEditLeftBTopWidth<HeightAnchorsakLeftakTopakRight TabOrder TextContentsNameEdit  TMemoContentsMemoLeftTop0WidthvHeightAnchorsakLeftakTopakRightakBottom Lines.StringsContentsMemo TabOrder    TPanel	SitePanelLeft Top Width�HeightaAlignalClient
BevelOuterbvNoneTabOrder
DesignSize�a  	TGroupBox
BasicGroupLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionSessionTabOrder 
DesignSize�  TLabelLabel1LeftTopEWidth=HeightCaption   &Värdnamn:FocusControlHostNameEdit  TLabelLabel2LeftTopEWidthFHeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlPortNumberEdit  TLabelUserNameLabelLeftToptWidth;HeightCaption   &Användarnamn:FocusControlUserNameEdit  TLabelPasswordLabelLeft� ToptWidth5HeightCaption   &Lösenord:FocusControlPasswordEdit  TLabelLabel22LeftTopWidthEHeightCaption&Filprotokoll:FocusControlTransferProtocolCombo  TLabel	FtpsLabelLeft� TopWidth<HeightCaption&Kryptering:FocusControl	FtpsCombo  TLabelWebDavsLabelLeft� TopWidth<HeightCaption&Kryptering:FocusControlWebDavsCombo  TPanelBasicS3PanelLeftTop� WidthvHeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
DesignSizev  	TCheckBoxS3CredentialsEnvCheck3LeftTopWidth� HeightAnchorsakLeftakTopakRight Caption'   &Inloggningsuppgifter från AWS-miljö:TabOrder OnClickS3CredentialsEnvCheck3Click  	TComboBoxS3ProfileComboLeft� Top WidthyHeightDropDownCountTabOrderTextS3ProfileComboOnChangeS3ProfileComboChange   TEditEncryptionViewLeft� Top(Width� HeightTabOrderOnChangeTransferProtocolComboChange  TEditTransferProtocolViewLeftTop(Width� HeightTabOrderOnChangeTransferProtocolComboChange  TEditHostNameEditLeftTopWWidth
HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderTextHostNameEditOnChange
DataChangeOnExitHostNameEditExit  TEditUserNameEditLeftTop� Width� Height	MaxLength� TabOrderTextUserNameEditOnChange
DataChange  TPasswordEditPasswordEditLeft� Top� Width� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextPasswordEditOnChange
DataChange  TUpDownEditPortNumberEditLeftTopWWidthfHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrderOnChangePortNumberEditChange  	TComboBoxTransferProtocolComboLeftTop(Width� HeightStylecsDropDownListTabOrder OnChangeTransferProtocolComboChangeItems.StringsSFTPSCPFTPWebDAV	Amazon S3   	TComboBox	FtpsComboLeft� Top(Width� HeightStylecsDropDownListTabOrderOnChangeEncryptionComboChangeItems.StringsIngen krypteringTLS/SSL Implicit encryptionXTLS/SSL Explicit encryptionX   	TComboBoxWebDavsComboLeft� Top(Width� HeightStylecsDropDownListTabOrderOnChangeEncryptionComboChangeItems.StringsNo encryptionXTLS/SSL Implicit encryptionX   TPanelBasicFtpPanelLeftTop� WidthvHeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder	 	TCheckBoxAnonymousLoginCheckLeftTop Width� HeightCaption&Anonym inloggningTabOrder OnClickAnonymousLoginCheckClick   TPanelBasicSshPanelLeftTop� Width�Height AnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder
  TButtonAdvancedButtonLeftTop� WidthlHeightActionSessionAdvancedActionAnchorsakRightakBottom StylebsSplitButtonTabOrderOnDropDownClickAdvancedButtonDropDownClick  TButton
SaveButtonLeftTop� WidthlHeightActionSaveSessionActionAnchorsakLeftakBottom StylebsSplitButtonTabOrderOnDropDownClickSaveButtonDropDownClick  TButtonEditCancelButtonLeftzTop� WidthPHeightActionEditCancelActionAnchorsakLeftakBottom TabOrderOnDropDownClickSaveButtonDropDownClick  TButton
EditButtonLeftTop� WidthlHeightActionEditSessionActionAnchorsakLeftakBottom TabOrderOnDropDownClickSaveButtonDropDownClick   	TGroupBox	NoteGroupLeftTopWidth�HeightNAnchorsakLeftakTopakRightakBottom Caption
AnteckningTabOrder
DesignSize�N  TMemoNoteMemoLeftTopWidthwHeight4TabStopAnchorsakLeftakTopakRightakBottom 
BevelInnerbvNone
BevelOuterbvNoneBorderStylebsNoneLines.StringsNoteMemo 
ScrollBars
ssVerticalTabOrder     TPanelButtonPanelLeft TopaWidth�Height"AlignalBottom
BevelOuterbvNoneTabOrderOnMouseDownPanelMouseDown
DesignSize�"  TButtonLoginButtonLeftqTopWidthlHeightActionLoginActionAnchorsakRightakBottom Default	ImagesActionImageListModalResultStylebsSplitButtonTabOrder OnDropDownClickLoginButtonDropDownClick  TButtonCloseButtonLeft� TopWidthPHeightAnchorsakRightakBottom Cancel	Caption   StängModalResultTabOrder  TButton
HelpButtonLeft9TopWidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick    TPanel
SitesPanelLeft Top Width�Height�AlignalClient
BevelOuterbvNoneTabOrder
DesignSize��  	TTreeViewSessionTreeLeftTopWidth�HeightVAnchorsakLeftakTopakRightakBottom DoubleBuffered	DragModedmAutomaticHideSelectionIndentParentDoubleBufferedParentShowHint	RowSelect	ShowHint	ShowRootSortTypestBothTabOrder OnChangeSessionTreeChange
OnChangingSessionTreeChangingOnCollapsedSessionTreeExpandedCollapsed	OnCompareSessionTreeCompareOnContextPopupSessionTreeContextPopupOnCustomDrawItemSessionTreeCustomDrawItem
OnDblClickSessionTreeDblClick
OnDragDropSessionTreeDragDropOnEditedSessionTreeEdited	OnEditingSessionTreeEditing	OnEndDragSessionTreeEndDragOnExitSessionTreeExitOnExpandingSessionTreeExpanding
OnExpandedSessionTreeExpandedCollapsed	OnKeyDownSessionTreeKeyDown
OnKeyPressSessionTreeKeyPressOnMouseDownSessionTreeMouseDownOnMouseMoveSessionTreeMouseMoveOnStartDragSessionTreeStartDrag  TButtonManageButtonLeftdTopdWidthlHeightAnchorsakRightakBottom Caption&HanteraTabOrderOnClickManageButtonClick  TButtonToolsMenuButtonLeftTopdWidthlHeightAnchorsakLeftakBottom Caption&VerktygTabOrderOnClickToolsMenuButtonClick  TPanelSitesIncrementalSearchPanelLeftTop5Width� HeightAnchorsakLeftakRightakBottom 
BevelOuterbvNone	PopupMenuSitesIncrementalSearchPopupMenuTabOrderOnContextPopup'SitesIncrementalSearchPanelContextPopup TStaticText!SitesIncrementalSearchBorderLabelLeft Top Width� HeightAlignalClientAutoSizeBorderStyle	sbsSingleTabOrder   TStaticTextSitesIncrementalSearchLabelLeftTopWidth� HeightCaptionSitesIncrementalSearchLabelShowAccelCharTabOrder    TPanelShowAgainPanelLeft Top�WidthiHeightAlignalBottom
BevelOuterbvNoneTabOrderOnMouseDownPanelMouseDown 	TCheckBoxShowAgainCheckLeftTop Width�HeightCaptionO   &Visa inloggningsdialogrutan vid start och när den sista sessionen är stängdChecked	State	cbCheckedTabOrder OnClickShowAgainCheckClick   TActionList
ActionListImagesActionImageListOnUpdateActionListUpdateLeft,Top TActionEditSessionActionCategorySessionsCaption	&Redigera	OnExecuteEditSessionActionExecute  TActionSaveAsSessionActionCategorySessionsCaption
&Spara somShortCutA�  	OnExecuteSaveAsSessionActionExecute  TActionSaveSessionActionCategorySessionsCaption	&Spara...	OnExecuteSaveSessionActionExecute  TActionDeleteSessionActionCategorySessionsCaptionTa &bort...
ImageIndex	OnExecuteDeleteSessionActionExecute  TActionImportSessionsActionCategorySessionsCaption&Importera...	OnExecuteImportSessionsActionExecute  TActionLoginActionCategorySessionCaptionLogga in
ImageIndex 	OnExecuteLoginActionExecute  TActionAboutActionCategoryOtherCaption&Om...	OnExecuteAboutActionExecute  TActionCleanUpActionCategoryOtherCaption&Rensa applikationsdata...	OnExecuteCleanUpActionExecute  TActionResetNewSessionActionCategorySessionsCaption   Å&terställ	OnExecuteResetNewSessionActionExecute  TActionSetDefaultSessionActionCategorySessionsCaption   Sä&tt som standard	OnExecuteSetDefaultSessionActionExecute  TActionDesktopIconActionCategorySessionsCaptionSkrivbords&ikon	OnExecuteDesktopIconActionExecute  TActionSendToHookActionCategorySessionsCaption"   Utforskarens 'Skicka till'-genväg	OnExecuteSendToHookActionExecute  TActionCheckForUpdatesActionTagCategoryOtherCaption   Sök efter &uppdateringar
ImageIndex?	OnExecuteCheckForUpdatesActionExecute  TActionRenameSessionActionCategorySessionsCaption	Byt &namn
ImageIndex	OnExecuteRenameSessionActionExecute  TActionNewSessionFolderActionCategorySessionsCaptionN&y katalog...
ImageIndex	OnExecuteNewSessionFolderActionExecute  TActionRunPageantActionCategoryOtherCaption   Kör &Pageant	OnExecuteRunPageantActionExecute  TActionRunPuttygenActionCategoryOtherCaption   Kör PuTTY&gen	OnExecuteRunPuttygenActionExecute  TActionImportActionCategoryOtherCaption'   Importera/Återställ &konfiguration...	OnExecuteImportActionExecute  TActionExportActionCategoryOtherCaption-   &Exportera/Säkerhetskopiera konfiguration...	OnExecuteExportActionExecute  TActionPreferencesActionCategoryOtherCaption   &Inställningar...	OnExecutePreferencesActionExecute  TActionEditCancelActionCategorySessionCaption&Avbryt	OnExecuteEditCancelActionExecute  TActionSessionAdvancedActionCategorySessionCaption&Avancerad...	OnExecuteSessionAdvancedActionExecute  TActionPreferencesLoggingActionCategoryOtherCaption&Loggning...	OnExecutePreferencesLoggingActionExecute  TActionCloneToNewSiteActionCategorySessionCaption&Klona till ny webbplats	OnExecuteCloneToNewSiteActionExecute  TActionPuttyActionCategorySessionCaption   Öppna i &PuTTY
ImageIndexSecondaryShortCuts.StringsShift+Ctrl+P ShortCutP@	OnExecutePuttyActionExecute  TActionPasteUrlActionCategorySessionsCaptionKlistra in sessions-&URLShortCutV@	OnExecutePasteUrlActionExecute  TActionGenerateUrlAction2CategorySessionsCaption&Skapa sessions-URL/kod...	OnExecuteGenerateUrlAction2Execute  TActionCopyParamRuleActionCategorySessionsCaption#   Överföringsinställnings&regel...	OnExecuteCopyParamRuleActionExecute  TActionSearchSiteNameStartOnlyActionCategoryOtherCaption$   Endast &början av webbplatsens namn	OnExecute$SearchSiteNameStartOnlyActionExecute  TActionSearchSiteNameActionCategoryOtherCaption&Varje del av webbplatsens namn	OnExecuteSearchSiteNameActionExecute  TActionSearchSiteActionCategoryOtherCaption   Alla &fält för webbplatsen	OnExecuteSearchSiteActionExecute  TActionSessionRawActionCategorySessionCaption   Redigera Raw-inställningar...	OnExecuteSessionAdvancedActionExecute  TActionSearchSiteStartActionCategoryOtherCaption&Hitta webbplatsSecondaryShortCuts.StringsAlt+F7F3 ShortCutF@	OnExecuteSearchSiteStartActionExecute   
TPopupMenuToolsPopupMenuLeft� TopM 	TMenuItemImport1ActionImportSessionsAction  	TMenuItemN3Caption-  	TMenuItemImportConfiguration1ActionImportAction  	TMenuItemExportConfiguration1ActionExportAction  	TMenuItemCleanup1ActionCleanUpAction  	TMenuItemN2Caption-  	TMenuItemPageant1ActionRunPageantAction  	TMenuItem	Puttygen1ActionRunPuttygenAction  	TMenuItemN1Caption-  	TMenuItemCheckForUpdates1ActionCheckForUpdatesAction  	TMenuItemN4Caption-  	TMenuItemPreferences1ActionPreferencesAction  	TMenuItemAbout1ActionAboutAction   TPngImageListSessionImageList	PngImages
BackgroundclWhiteNameUnusedPngImage.Data
b   �PNG

   IHDR         ��h6   tRNS �   ���/�   IDATx�c����8�aT���  �E�/UY"    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
k  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:04+01:00" xmp:MetadataDate="2022-09-01T11:08:04+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:90551216-ab82-2c46-b9c8-b8ddacc04ba4" xmpMM:DocumentID="adobe:docid:photoshop:c10ce5f3-4426-6940-933a-9d2fd6bcda2d" xmpMM:OriginalDocumentID="xmp.did:4442d8a0-33db-2a47-9031-55ffc0f53f64"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:4442d8a0-33db-2a47-9031-55ffc0f53f64" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:90551216-ab82-2c46-b9c8-b8ddacc04ba4" stEvt:when="2022-09-01T11:08:04+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>rTb  HIDATx�c���?%�d@�)/���+���? �(| �B�Ŕ���p:{&�������?0���1�����3�L`������[0ÿ��4��0����93� hl����-�������1,�3a@mC����x5�]t�۵�K�APY���KT����|}�ʥ�V��������|���֮\�0�����.�x^��a����׮D�[P��cQ����͉[7�E��]��߿�"��?h��������j���p�&����yFj"�X�j��-;���޾󅄅�t��#Q�{�c�a;�n�n Ź�  ?@��y�ؕ    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:08+01:00" xmp:MetadataDate="2022-09-01T11:06:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5f0285a2-1a20-234b-9a43-8da79e79cb07" xmpMM:DocumentID="adobe:docid:photoshop:9a4cfe93-5052-9246-bf53-fd91397c86e1" xmpMM:OriginalDocumentID="xmp.did:ed00465a-0d10-4b4e-a04b-d555174bc285"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ed00465a-0d10-4b4e-a04b-d555174bc285" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5f0285a2-1a20-234b-9a43-8da79e79cb07" stEvt:when="2022-09-01T11:06:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Z��  �IDATxڭS9KQ���l�V�PW#*Z��I�Bk� Z��o�j����^�Q�� o���&;Ƹ� t�ͼ���73���3��V���T c�q)p5�;�U%�46�=���vI'��C���T�����?URq�Ͽ���I[Q�8G����X�*A�N8��Y���۲�B�R��W��`����+`j@\KZ�,$y���~�:�����3� `;p����(���iTF]k��JГ���8��ȼa������S	vDdj�^x�����$l��iSϪ�IS�t��{�|�����֮�<լqr��	)p��7;K�Q�؞�Z�8������j�v����Cy�l�ai"==L��Q[����)����Q^�~�@�F����_�� &M?�ZP    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:06+01:00" xmp:MetadataDate="2022-09-01T11:02:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:72f8666d-2ee5-344b-aa1d-a1c6ea8cd32b" xmpMM:DocumentID="adobe:docid:photoshop:cba89235-7918-cb4d-9b5c-ca3e0435cf2a" xmpMM:OriginalDocumentID="xmp.did:7bb19fbd-fb7b-5f47-87b8-73ea5303e6e4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7bb19fbd-fb7b-5f47-87b8-73ea5303e6e4" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:72f8666d-2ee5-344b-aa1d-a1c6ea8cd32b" stEvt:when="2022-09-01T11:02:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��t�  mIDATx�c���?%���N!Y&� �?_ZO�:�����F�Ō�wK�2�Pe���=�!ʀ_����P���?�=�r��;� �1~ކ� fNqf.i �� ���������\N�y���f���K�j�$3��6���oH�����������X�6��ݮ����a`��*�����{������4�����fje�91��Z���:L��!
�h���r��4��]�WJ��5L���M3�fuy�d�~$A(.z���)� � �6��P��"�g�8T3���5�h���NP��j����4���Q5��6�7Ԁ+��32��d~$:20ܒ{
�+��fg }6�e>M    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:10+01:00" xmp:MetadataDate="2022-09-01T11:08:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:1f1a0273-57ab-fe41-ae28-870eeaf05b00" xmpMM:DocumentID="adobe:docid:photoshop:81d5b2de-52b0-0544-9841-c4936f1aa521" xmpMM:OriginalDocumentID="xmp.did:878c169a-9444-1047-bff4-907f81185561"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:878c169a-9444-1047-bff4-907f81185561" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:1f1a0273-57ab-fe41-ae28-870eeaf05b00" stEvt:when="2022-09-01T11:08:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>X�S�   �IDATx�c���?%�Q��-�L`T[{�2�͜���ۋ,�[�n�����U��Y�p����d$D3�~v��MACAJJ4ëo�y�q��a��!�A~�9� �l���m&\H`�>�"�j [�^ �1|�������lc���r&��n�.�eHAzR�����Eq� �- v\P"åU�,����h���&+!=��J)�,�P�Hiv B����    IEND�B`� 
BackgroundclWindowNameWorkspace closed (unused)PngImage.Data
b   �PNG

   IHDR         ��h6   tRNS �   ���/�   IDATx�c����8�aT���  �E�/UY"    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
-  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:07+01:00" xmp:MetadataDate="2022-09-01T11:08:07+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c152f702-baba-cc4c-a6b8-23ee1a3c60a0" xmpMM:DocumentID="adobe:docid:photoshop:386766ec-32ad-9948-9e34-76bdeb9fddb2" xmpMM:OriginalDocumentID="xmp.did:7164580e-2ba8-3146-8f84-f140a4cc7694"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7164580e-2ba8-3146-8f84-f140a4cc7694" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c152f702-baba-cc4c-a6b8-23ee1a3c60a0" stEvt:when="2022-09-01T11:08:07+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  
IDATx�c���?###!0s��<F&��g~�6����3��0��߿����� ����QPP`���a�y��۷o_L��'	7��g�����P���/�߿�3�|y�,�͠,#ɰ��5�;'0�+kI|���l@kG���n��~�����5���[̬�L@��C���^]�j-�E@������4�t����b;���/w��Y�l��� ^�7��2�;p���*��6���������A��s�0�@����ǰj�:�a��2����i���%
j�C��3���b����?�+6m���������K`J+j��p��kBvI:�}+eI��o>1|~��A^V����w>~��JOY6�����.�x/�p.0 �3���p�+�%�3���`��0 �����$���ߨ|�ۓ�lX�O�����+�)!��80 _�ܶQn ��<c��� :#5gZ�j��-;�߽}�	��@F�p����Ͷ�[7b7�@� ���ն�"    IEND�B`� 
BackgroundclWindowName Open new session closed (unused)PngImage.Data
r   �PNG

   IHDR         ��h6   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?)�qTè�� ��/�Ǭ�Y    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
D  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:01+01:00" xmp:MetadataDate="2022-09-01T11:08:01+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0a7dbdf9-638c-2a4c-871c-bf60320321c2" xmpMM:DocumentID="adobe:docid:photoshop:81b209e4-a2e5-1749-ba81-14162fdaf5d7" xmpMM:OriginalDocumentID="xmp.did:dbb80521-31b4-424d-a0fd-57346150a394"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:dbb80521-31b4-424d-a0fd-57346150a394" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0a7dbdf9-638c-2a4c-871c-bf60320321c2" stEvt:when="2022-09-01T11:08:01+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�͇�  !IDATx�c���?%�d@�)/���+���? �(| �B�Ŕ���p:{&�//- �֌��S&0�h���_]YB�)�9sfLA���񿾶�h�3̙�0����sc��ħ0,Y0a@eM�������gX�t!Ҋ��ݝ-DͰv�R��%��{;�6�?(�a�ڕrJ�O��C��~�[7�E �����AN8���[����߫[7��`dd�jӌ����<#5C,`5`��`�wo߂�B��`:�ǃ�(ܽ��氝[7b7�@� �v��t]��    IEND�B`�  Left,Top�   
TPopupMenuSaveDropDownMenuLeftTop 	TMenuItemSaveSessionMenuItemActionSaveSessionActionDefault	  	TMenuItemSaveAsSessionMenuItemActionSaveAsSessionAction  	TMenuItemN7Caption-  	TMenuItemSetdefaults1ActionSetDefaultSessionAction   
TPopupMenuManageSitePopupMenuImagesActionImageListLeft�Top 	TMenuItem
Shellicon1Caption	WebbplatsEnabledVisible  	TMenuItemSiteLoginMenuItemActionLoginActionDefault	  	TMenuItemOpeninPuTTY2ActionPuttyAction  	TMenuItemN10Caption-  	TMenuItemEdit1ActionEditSessionAction  	TMenuItemDelete1ActionDeleteSessionAction  	TMenuItemRename1ActionRenameSessionAction  	TMenuItemSiteClonetoNewSiteMenuItemActionCloneToNewSiteAction  	TMenuItemGenerateSessionURL1ActionGenerateUrlAction2  	TMenuItemN5Caption-  	TMenuItemSetdefaults2ActionSetDefaultSessionAction  	TMenuItemN6Caption-  	TMenuItem
Newfolder1ActionNewSessionFolderAction  	TMenuItem
Shellicon2CaptionIkon webbplatsEnabledVisible  	TMenuItemDesktopIcon2ActionDesktopIconAction  	TMenuItemExplorersSendToShortcut2ActionSendToHookAction  	TMenuItemSearch1Caption   SökEnabledVisible  	TMenuItem	FindSite1ActionSearchSiteStartAction  	TMenuItemSearchOptions1Caption
Alternativ 	TMenuItemSearchSiteNameStartOnly1ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemSearchSiteName1ActionSearchSiteNameAction	RadioItem	  	TMenuItemSearchSite1ActionSearchSiteAction	RadioItem	    
TPopupMenuManageFolderPopupMenuImagesActionImageListLeft�TopM 	TMenuItem	MenuItem1CaptionWebbplatskatalogEnabledVisible  	TMenuItemLogin5ActionLoginActionDefault	  	TMenuItemOpeninPuTTY4ActionPuttyAction  	TMenuItemN11Caption-  	TMenuItem	MenuItem3ActionDeleteSessionAction  	TMenuItem	MenuItem4ActionRenameSessionAction  	TMenuItem	MenuItem5Caption-  	TMenuItem	MenuItem6ActionNewSessionFolderAction  	TMenuItem	MenuItem7CaptionIkon webbplatskatalogEnabledVisible  	TMenuItem	MenuItem8ActionDesktopIconAction  	TMenuItemSearch3Caption   SökEnabledVisible  	TMenuItem	FindSite3ActionSearchSiteStartAction  	TMenuItemSearchOptions3Caption
Alternativ 	TMenuItemBeginningofSiteNameOnly2ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemAnyPartofSiteName2ActionSearchSiteNameAction	RadioItem	  	TMenuItemAllMajorSiteFields2ActionSearchSiteAction	RadioItem	    
TPopupMenuManageNewSitePopupMenuImagesActionImageListLeft� Top�  	TMenuItem
MenuItem12CaptionNy webbplatsEnabledVisible  	TMenuItemLogin2ActionLoginActionDefault	  	TMenuItemOpeninPuTTY3ActionPuttyAction  	TMenuItemN8Caption-  	TMenuItem
MenuItem13ActionSaveAsSessionAction  	TMenuItemReset1ActionResetNewSessionAction  	TMenuItemPaste1ActionPasteUrlAction  	TMenuItemGenerateSessionURL2ActionGenerateUrlAction2  	TMenuItem
MenuItem21Caption-  	TMenuItem
MenuItem22ActionSetDefaultSessionAction  	TMenuItem
MenuItem16Caption-  	TMenuItem
MenuItem17ActionNewSessionFolderAction  	TMenuItemSearch2Caption   SökEnabledVisible  	TMenuItem	FindSite2ActionSearchSiteStartAction  	TMenuItemSearchOptions2Caption
Alternativ 	TMenuItemBeginningofSiteNameOnly1ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemAnyPartofSiteName1ActionSearchSiteNameAction	RadioItem	  	TMenuItemAllMajorSiteFields1ActionSearchSiteAction	RadioItem	    
TPopupMenuManageWorkspacePopupMenuImagesActionImageListLeft�Top�  	TMenuItem	MenuItem2Caption	ArbetsytaEnabledVisible  	TMenuItemLogin3ActionLoginActionDefault	  	TMenuItemN9Caption-  	TMenuItem
MenuItem10ActionDeleteSessionAction  	TMenuItem
MenuItem11ActionRenameSessionAction  	TMenuItem
MenuItem18CaptionIkon arbetsytaEnabledVisible  	TMenuItem
MenuItem19ActionDesktopIconAction  	TMenuItemSearch4Caption   SökEnabledVisible  	TMenuItem	FindSite4ActionSearchSiteStartAction  	TMenuItemSearchOptions4Caption
Alternativ 	TMenuItemBeginningofSiteNameOnly3ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItemAnyPartofSiteName3ActionSearchSiteNameAction	RadioItem	  	TMenuItemAllMajorSiteFields3ActionSearchSiteAction	RadioItem	    
TPopupMenuSessionAdvancedPopupMenuLeft� Top 	TMenuItemSession1CaptionSessionEnabledVisible  	TMenuItem	MenuItem9ActionSessionAdvancedActionDefault	  	TMenuItemEditRawSettings1ActionSessionRawAction  	TMenuItemTransferSettingsRule1ActionCopyParamRuleAction  	TMenuItem
MenuItem14Caption   Globala inställningarEnabledVisible  	TMenuItemPreferencesLoggingAction1ActionPreferencesLoggingAction   TPngImageListActionImageList	PngImages
BackgroundclWindowNameLoginPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:05+01:00" xmp:MetadataDate="2022-09-01T11:06:05+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f2062452-6d8e-0d48-bb77-752c4ec26b5a" xmpMM:DocumentID="adobe:docid:photoshop:a9199e92-8997-0442-b578-638372c4c5c1" xmpMM:OriginalDocumentID="xmp.did:ba568a23-305e-1045-9542-b55c9f2c5fde"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ba568a23-305e-1045-9542-b55c9f2c5fde" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f2062452-6d8e-0d48-bb77-752c4ec26b5a" stEvt:when="2022-09-01T11:06:05+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  �IDATxڥ��/A����U�zs�
Q�.����,� qt��(�&�"8xU��MۭnI<v�iZ:A"�m�;��o>3��K(�H$H�3����kd�u���`&�f6h I,]�j�}�����I�b@8iJ��H�<�~
����*� Ӥ�s��#V=S_���a��� �wu�� �^����^ܿ�`_v�mc�)��	W� �i�Y��_8�т���	<�2�-�(�f�� j5����I�v5�}�˭
�$<�@z���f�o�ˀ6���"P��~;���it�Z���K��7�����`�� �+U^Еg�>5ʛ��k��q��ҡ�]�r. �
�t�G �{*�F�+�
��$�.D�\�5�Y����~��|/�mU"t) iejlf���'�w`��%����sZ�B����	�t�r��    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
V  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:11+01:00" xmp:MetadataDate="2022-09-01T10:57:11+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0832a1ea-198f-ec43-9943-930a416eb7c8" xmpMM:DocumentID="adobe:docid:photoshop:55fb95e1-5c0b-8a4f-a24c-51622779ce43" xmpMM:OriginalDocumentID="xmp.did:5773b47b-d28d-2f45-8cce-bd07d1224e92"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5773b47b-d28d-2f45-8cce-bd07d1224e92" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0832a1ea-198f-ec43-9943-930a416eb7c8" stEvt:when="2022-09-01T10:57:11+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  3IDATxڅ�_HSQǿgӭ�Y$��bO����^"���!�P4�ПV�X�-���H2��cA�b2� ��RQ�䋤"�����v�=�s�Vʽt�ǹ���~��~���
/k�V���F)�{�[T�~%f�[�!6�����iv�'v��V=�{\�{MSO`
��b�'�XC���@4]�  n�zh����)�MO \B�����>�S�5>2�g��`eN�ٞ�f/���/?��C��p�����,�Սa_m���ӽԌ���`_T��=��a�d�X��e�,� �
5�Aۢs�j�Rd.b���]����t�c��@ͺ��:���?�����re��ɇ���\@���q��	� Mf�u�����9�*7"�Z��<d���W�X,BL�|rh�W
6UT����&	"��t�Qg���9��FK���V��u���@2�\5�ї�+����y&g]GiV�x�i����2D4Q-�|��p��{��#ܒ��j���}w"{��"��F�6�6z�1�z=gM/�!``8"���qð�hl>Ό6��2{� x�Z�"J�j    IEND�B`� 
BackgroundclWindowNameRename 2PngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:13+01:00" xmp:MetadataDate="2022-09-01T11:08:13+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ece3c1d3-e8ce-fc40-8183-104e6cbbf44f" xmpMM:DocumentID="adobe:docid:photoshop:8cb8788e-c0cc-1b42-8433-1838e2f16f65" xmpMM:OriginalDocumentID="xmp.did:8d0f831c-d906-c442-ac82-73cfc3e57db7"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8d0f831c-d906-c442-ac82-73cfc3e57db7" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ece3c1d3-e8ce-fc40-8183-104e6cbbf44f" stEvt:when="2022-09-01T11:08:13+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>w�e�  mIDATx�cd �IS����'ݏ�>d2�����\�G�������ߏ�d���,�f��=�xZ�ǄL~�g7=I2��q���LR�W�
�={��_h�/�|?b#������__�~�p��������D������x���蔟9ln/��ĉ2��1� ����������ogڎ>7oh`�G���k�s\����������e����L��������������~Ndsy^�,�8m����4s�gRZ� ����O&�Տ~�cc�0 3-	�6�3��d�d����?��Q�E~��y���;�/����;e�8Q���5���K;#�����"L�pb��o_>28�g�`Hp�� A۽ cOy/    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:50:59+01:00" xmp:MetadataDate="2022-09-01T10:50:59+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c52f6a03-faa9-0a4d-bab9-6c89b0f5b88a" xmpMM:DocumentID="adobe:docid:photoshop:540cb7cd-9414-c44b-8739-5ac78f6cc1ae" xmpMM:OriginalDocumentID="xmp.did:01e6ad1a-5a6e-2145-8135-0dca66c44d55"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:01e6ad1a-5a6e-2145-8135-0dca66c44d55" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c52f6a03-faa9-0a4d-bab9-6c89b0f5b88a" stEvt:when="2022-09-01T10:50:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��^  yIDATxڭ��K�@�_�ڦź���U��:�n�.
��������A�NF\�;�ME�mM�����]���V
�7�}>���;��`�R�M�~�����f�>̕�����vF�Njet���U�*	��%�}��-#*p:��@����U�o��PM@�!s>:F�&���c���ՊmIEQ�u^WT�$�H�Zͮ�q7�׮��
D		 ��@b|=��,�~>2j�`C+�g� ��^����	�;�����v_2R���bMC�D�q|b^�1r�`	�vf���̵BFO�(�;<~����%������H��%�ǧ�&�`e���+	�K���J�m�+E�AI,��p]:Y���Wy������+K�|�6    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
6  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:51:04+01:00" xmp:MetadataDate="2022-09-01T10:51:04+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d01c1147-26b2-2d4f-ab0a-36111a1c0ea2" xmpMM:DocumentID="adobe:docid:photoshop:54c5e437-fdec-1f47-a95f-b644f5e3c30d" xmpMM:OriginalDocumentID="xmp.did:03e4f68b-4129-8f4c-8a95-6ad9e03db62b"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:03e4f68b-4129-8f4c-8a95-6ad9e03db62b" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d01c1147-26b2-2d4f-ab0a-36111a1c0ea2" stEvt:when="2022-09-01T10:51:04+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>j�H�  IDATxڕ�OhAƿצ�h���d�"��ؠ ��V0B�S�
-(�֐���ă�@�"JUP�R���A+���VhS�Jk$��v7�;�t�lk%>�c����7�%�1�޻�P\/XF�DB�}Oj�����@p{.Ț��\�4�
�_�>���?���_�;�m0���$�"R����hRQ�[_O����Y:��1��gK��"��v�����۳�{�H�&F)%��%������Q�>�^`%�\�؏$l_' �2c����P����a��M��F8��+���Al	��A����}�ˁ��0��	L�]L^�{@�젠�����k��".�ю�ǎ����ёgPU#�J�'��m|G4i�`:��;�j���I4��C_�cn^���$�����D�C23��ȁ>p�J�Nv��{� "�d��ԘU�p]T�kDmF�?�sv�h�w������Ru�B�@�G�8���^���Gp�Xٳ'������ݙ�M1E���I����������N-���u���]�~�9    IEND�B`� 
BackgroundclWindowNameOpen Workspace (reduced alpha)PngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06+01:00" xmp:MetadataDate="2022-09-01T11:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:dc9f4636-e72f-b241-8feb-bff3a506734e" xmpMM:DocumentID="adobe:docid:photoshop:71703c92-58e0-3b43-9912-7fdd1f3e4a03" xmpMM:OriginalDocumentID="xmp.did:e297fbb5-2a1f-894f-b2d5-a1cf3d391ad9"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e297fbb5-2a1f-894f-b2d5-a1cf3d391ad9" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:dc9f4636-e72f-b241-8feb-bff3a506734e" stEvt:when="2022-09-01T11:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>WpT�  �IDATx�cd@�ۯ�g \��ddD�6s�oo/���n�����cV�_{$�0�gԆI̹�̐��W���0��Ɂ>kCVz2#��R(N�p�_�Ai�3�������c#Q�X 1梹 �~ERQ�`�Rŕ��?v �1�1Ê�`JV;3��w10�~���Ȃ5��|������̂lJ�@!�0������k` <f���@�����Ci6Ὄ��I���f����OU���_��)F�#�%��H��Q�AFӍA@X��'X!����f��n���;ϙ�XXX���k�f�������r�����1��d`q�O��b�����-s�'���� i��6�w0�������j���<2�:8mC�\�w(���5��+��U5g��`�~"�������_��no�1��.����������LJ-'�Z�����{� ��[
lݾ�    IEND�B`� 
BackgroundclWindowName"Open saved session (reduced alpha)PngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:57:55+01:00" xmp:ModifyDate="2022-09-01T10:52:51+01:00" xmp:MetadataDate="2022-09-01T10:52:51+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9c7001f2-79d1-a948-bd21-bd3ed0bf3afc" xmpMM:DocumentID="adobe:docid:photoshop:08761404-3b30-e442-91bb-25734b9383d6" xmpMM:OriginalDocumentID="xmp.did:08b74781-ce3b-114b-a894-5582f1fdf500"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:08b74781-ce3b-114b-a894-5582f1fdf500" stEvt:when="2022-06-27T15:57:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9c7001f2-79d1-a948-bd21-bd3ed0bf3afc" stEvt:when="2022-09-01T10:52:51+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>F  �IDATxڍ�MHTQ���y3���2!�Ҩȅ(8�d�l7A$Em#re���FQ(Aٺ6~�A�h�BrӠ�>6�6JaM꼏����7��!/��?�q��s��ʬ���B�:)��T�R�Q9���Ou_�0S�[��=;�IL��#K`j�	,��x��Ùxo.Y� ����
�V���-s�}߁���ƬI��%_zT`ﳫ�n��ś�1"Ӑji��8
K<�o`�QT;�p�n���YtʀH��߫��k��1�N��k>׎ 쟀�Gl�	5�����Jh��ۡ���e���J��>�Eg/���آԬ��SQ�7�Qm����?�t;mL��5@��mh�V�`�~ rL�S�c5�Ϝ�oIm�w|ڴ�*�����ie��S���3=e�y��c���{��Y����DK�jE���ez�]k�)��874�C�6�{ay��2l����A�?�U�He8��.�Z�][=��̼o���ұ2H�/    IEND�B`�  Left)Top�   
TPopupMenuLoginDropDownMenuImagesActionImageListLeftTopM 	TMenuItemLogin1ActionLoginActionDefault	  	TMenuItemOpeninPuTTY1ActionPuttyAction   TPngImageListSessionImageList120HeightWidth	PngImages
BackgroundclWindowNameUnusedPngImage.Data
v   �PNG

   IHDR         �Z   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?��qT��Qͣ�V3 O�;ه>�    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:05+01:00" xmp:MetadataDate="2022-09-01T11:08:05+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d5ba6480-fce4-8340-bab0-dc63bbeea569" xmpMM:DocumentID="adobe:docid:photoshop:c6ddd208-eea0-fd4e-8f53-c64a5a5f8aea" xmpMM:OriginalDocumentID="xmp.did:00eaba8c-2121-a841-8bd1-5acdf139ff5e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:00eaba8c-2121-a841-8bd1-5acdf139ff5e" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d5ba6480-fce4-8340-bab0-dc63bbeea569" stEvt:when="2022-09-01T11:08:05+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�u�Y  �IDATx�c���?5#����S����O�@�/�����PLCő�_T��)z��v�M���͟����A����9�82��ϕ�ӧL`������[ �_AV�}u!ì��t��������!�^��3̝5a`ck���.!�^%`�E���1,�;a`]S��-�a���!��n7�0,Y0a`u]���Α���7��r�9�a���+���os��Ԁ�uh��ܚ��j�"���5�w8�`�տ\��oOgX�r)������;�Ȉ���T�kV �+*���!�V�^ƴ���d���W#��/��FhY�/�l�";���Y�öM�fd�����:�@�yU������7wlݠ7���g�1s�xq����S!���j��-;���{�..$,g�x0�e .@�����ܹu#n�	�n  t���pR��    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:09+01:00" xmp:MetadataDate="2022-09-01T11:06:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c9283f14-3d59-ec42-94c8-a53f7ac56617" xmpMM:DocumentID="adobe:docid:photoshop:39bb9190-aaa7-5f45-8ad3-4816d448e4c3" xmpMM:OriginalDocumentID="xmp.did:8f445be8-9da7-1a46-99ef-30686812fd01"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8f445be8-9da7-1a46-99ef-30686812fd01" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c9283f14-3d59-ec42-94c8-a53f7ac56617" stEvt:when="2022-09-01T11:06:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��Q5  �IDATx��MOA�����R���z��F�Ҙ� B?��iL<y ��K4�WCԛH0��Xhm�����<l���mnN��ϼ<��?��#"\fc�)��ap��	P�=�3�//|k+�&	��M���Z�Rb���7��b
��Ѱ�j���"zo'��r��=+�I�A>(S�B�9����:�KV./��F]�:��j�Ջ�� ֑c���A��S%��q��_��?�u`I�
�igAE.�'�A��r��y	<~�oʼ���[��������f�eF%���UY7v�8�d����v�A�L��ԇ�F$��&F'4��#ݸ�|L��-��l`�|�N~}*��5�
�~�)�E����_0ތ��_��ΒV��
���9�~n��U��q<2�sOWG�G��xz�-��g����g���I�.��]������~ReI���{���a�1�D�Ѷ���V���������˫�ҵ�v=���ul�L.��l�pP�q�r{    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:07+01:00" xmp:MetadataDate="2022-09-01T11:02:07+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:97d12c2e-ed65-a447-958b-fe256ac98664" xmpMM:DocumentID="adobe:docid:photoshop:469e9482-7664-3f42-92cf-ba17ffa1700a" xmpMM:OriginalDocumentID="xmp.did:62777e29-adc1-d44f-acc9-9c4ebedb8b10"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:62777e29-adc1-d44f-acc9-9c4ebedb8b10" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:97d12c2e-ed65-a447-958b-fe256ac98664" stEvt:when="2022-09-01T11:02:07+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>6�L  �IDATx�c���?5��0��.aY&d	����|u����!C�6���@!!L�S�ܞ�l��=��������Ny�wٝ_�#�@&qFi ����Q��_~e��̃b����Y9� ���Ҍ,���<r�C�����P�����A��������������] j;�п��g`������@�?�f�ߟ63!��T��S�/�����V��/B!>�pV�[�>Z%�_�8��M.>̥�N�h����k���.O�����ho���2��x�	������:�a�������*v�<��Q�����$~�j8��~c�&���� m*��L������e��0�0���|�R�:#��O@�GB%: �tK6�i��� ����0    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:11+01:00" xmp:MetadataDate="2022-09-01T11:08:11+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:98124c18-191b-b244-a7d5-4a004b509180" xmpMM:DocumentID="adobe:docid:photoshop:ecaf6699-1198-a345-be71-69e684951c09" xmpMM:OriginalDocumentID="xmp.did:d562b312-1a72-7040-b236-86d61f7228ca"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d562b312-1a72-7040-b236-86d61f7228ca" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:98124c18-191b-b244-a7d5-4a004b509180" stEvt:when="2022-09-01T11:08:11+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���   �IDATx�c���?5����T5�Q{�u����2u�6s�oo/���n��@HL��̴$�
�Ϛ�@HL��[v,`A�Cp���_���4A0 ��f ���e|ށ�{�4����4qy�@�{�w`���5q�f ./#H_/KJKTLx��)qy�X ��T1
�^bS�@ ��M��d6    IEND�B`� 
BackgroundclWindowNameWorkspace closed (unused)PngImage.Data
v   �PNG

   IHDR         �Z   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?��qT��Qͣ�V3 O�;ه>�    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:08+01:00" xmp:MetadataDate="2022-09-01T11:08:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ea9c212b-5fdb-6c42-b036-564a59974ad5" xmpMM:DocumentID="adobe:docid:photoshop:efebda47-97d3-994f-8c20-c0875567e635" xmpMM:OriginalDocumentID="xmp.did:38a4f023-e13c-e642-acc7-db653a64d539"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:38a4f023-e13c-e642-acc7-db653a64d539" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ea9c212b-5fdb-6c42-b036-564a59974ad5" stEvt:when="2022-09-01T11:08:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  �IDATxڭ�mHSQ�����eiP2��C�!�#|)z������5cYaY�aK*���з0��m�e�)A�^4́X���R9w�9����nmS1<��<���}^�s8�8��bV]C�&�B�+,���|��g���SJ׋��&T<��s�%j��cc0�ɌA������w6���:֔�D�@����|g���e38qh?M�h���������˚S�A�DO�D?�`~T@f��
��jţ�VpD�J��`&	x��6kݕ္��v�i���u�);�#0p9�>��B%p_�G:b��J�k7n�����������u �	񈉌p֒9j-�W�7���N�/+*o����>��Q�{��4�mf�d��7>6�	$^�;�Z�WT2S��T���$�Cα,'��]7<1bZ�,-��:���v�+�2���o �_F�6<[�"���%ld6�H���%�WXgR�o�����rE�B��!x5���?H�� �m+*�#�K�XWR�߆�#d��S㕘�)�?&^#͸�ua
�^O%����yb�ۙ������߉C���lp_l���L-��#^c�)a�Ni~�_N��6�X�;7H�(=���3,]rF����%J�����lmAނϒ_���S�L�����CCe;}�s�Ew��,�2��\ʵ������2 ���    IEND�B`� 
BackgroundclWindowName Open new session closed (unused)PngImage.Data
v   �PNG

   IHDR         �Z   sRGB ���   	pHYs  �  ��o�d   IDATx�c���?��qT��Qͣ�V3 O�;ه>�    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:02+01:00" xmp:MetadataDate="2022-09-01T11:08:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:960457fd-f233-b043-b30c-0ea7b39f277e" xmpMM:DocumentID="adobe:docid:photoshop:39028b26-ea30-3342-91b5-08c919050f10" xmpMM:OriginalDocumentID="xmp.did:93983595-bf6b-0449-a695-4a66d970cb9e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:93983595-bf6b-0449-a695-4a66d970cb9e" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:960457fd-f233-b043-b30c-0ea7b39f277e" stEvt:when="2022-09-01T11:08:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>˞��  rIDATxڭ��J�A ��W�^�n�9�)�Ȑ$I�V-�L���45MQ3K%iߵŰ7�����������L�?�����3g0 �v����!���HLAl��Z�����B��=��vS0K��l�բވҩ�`(�u�\�-�lz���P\�5npv~	�����q�s��-*�3t����8�A��:.��t� ���U�itvt�@�����T�&���!-6D�~nP��@7'4Y��nq�r�8*]�3�`�B2�����C��3�2�UrB��kd�F�~8����-uz��CA�m^�����J��KA���s2����sɍ�_�%X|�P�Z��2�`.P*����	>���vF��/�8����    IEND�B`�  Left� Top�   TPngImageListActionImageList120HeightWidth	PngImages
BackgroundclWindowNameLoginPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:06+01:00" xmp:MetadataDate="2022-09-01T11:06:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:3ad8c394-c1ef-2b4f-a5d6-629ca2484f69" xmpMM:DocumentID="adobe:docid:photoshop:43507e1f-292a-6440-8cfb-11aa6d58b35b" xmpMM:OriginalDocumentID="xmp.did:e5f48a6f-60a5-c94f-8cfb-489c78fabfc0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e5f48a6f-60a5-c94f-8cfb-489c78fabfc0" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:3ad8c394-c1ef-2b4f-a5d6-629ca2484f69" stEvt:when="2022-09-01T11:06:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>+K��  uIDATxڭ��ORa��A�$��h��-��j�Q�[fu��*/�Rֵ�ռ���es�F��VʹF[4�/����"�� �����}��y���{�� ��bb��.��1b3�B��l�&��Ba_OxY���,����(����2Ϥ�b��)@{JF�l��K�Z����
�)��6���ザsao��Ʌ��r8&o��ߓ����K���ԳM�=ܐ5Z��V}��9;^�"��k��S�j�9m+���X��2�8m��ex�Q��G�J��������^Ɩ\b�Dc�ލ�~�@�$V��&�"-���uN>y�7ۍ��;R����jƆ�o4X�ì���:놿[ ���-]t��	Ί���s0�^Õ��a\ ����8m��0Vq`��-�+ ��������Ƴ	qˤǚ�8B��9���v�U���]�?��ȓH%?ik}v�$��(K���,07�֠	������m�P��t	8#�c��('5���4"��Z7���_6,��#)���M�0�3w�Ҩ���ӊ��,{(0�0'5�)`*��B�����h�|�����ݕE��f�����&���	9�@�`7S�`[�v+�}���E��    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:12+01:00" xmp:MetadataDate="2022-09-01T10:57:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:1f526019-6579-9349-b850-cca8486a5703" xmpMM:DocumentID="adobe:docid:photoshop:605cf25d-e29b-9d45-8ff3-e3c241e40fa7" xmpMM:OriginalDocumentID="xmp.did:9d390167-571b-8849-b77a-dc84de202c61"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:9d390167-571b-8849-b77a-dc84de202c61" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:1f526019-6579-9349-b850-cca8486a5703" stEvt:when="2022-09-01T10:57:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  �IDATxڕ�mHSQ��g�cKjf�!�1��!�`,��D"bFI%$*�,X���4C2��H􃐥�iH !�� �L�S$�%Y���r:wӵ9w�Ͻ��s���y��(\������K�$����.��o�QV�ܡ�S3!�%OHkO��Ko�"����v%!�� ����F��Xr�}д���7*��䬀L�ߡVk� R[�p�}�)-����
�{2ۗ����-�Ѕ��4s�%6O�묊䉇��k&3}���v�L��1l�V8l�H���Gl@�I���W�Mt4�4,��a�PqZ���|r�-��ց��� JjDi��w��z5���A�y}�Gϯ���>>� J���(긛�i���d��bu"~��w3�@m���jt����_Ā&�Ԡ�+D�1�v�l	��#X�i|��*��fjȱW�a�뚑��d)�,������1r[���lT�!�`hgt�j��I�fc^8�m��H�T����� h��%Qm���?��j8�a���@o�_��F�٠s��.��"��������A�	�����R7RRZN_�8X.O���Ce�=�)@�R<
?����<jtwv���AÅ �^��#�[@����fAXk��F_wgh��+�?��;D?��t�������c�s4����`=�		�����JT������?��z�����g���LIϠ�}识���&/پ`�K    IEND�B`� 
BackgroundclWindowNameRename 2PngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:14+01:00" xmp:MetadataDate="2022-09-01T11:08:14+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0f5181e5-1423-9340-922b-d3c5ac93e227" xmpMM:DocumentID="adobe:docid:photoshop:875c291a-6310-d940-8f09-f96d889da58b" xmpMM:OriginalDocumentID="xmp.did:fde8fd27-e4c0-074b-a37b-670b399d123d"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:fde8fd27-e4c0-074b-a37b-670b399d123d" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0f5181e5-1423-9340-922b-d3c5ac93e227" stEvt:when="2022-09-01T11:08:14+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��7  �IDATx�c���?###��M��������4Ef��Ō��r��/�??|f���;e~�t��ۖ�}ߎ�d ����\��p)J�Mu��W��ʾ߷��ʶO?��V%�������ar��U�����&�^+�NH�'����-���<���w ~��z��ǲ$������b�nr�ߟ�����_��on�e������h����iaw}^�'���Gl�������;ذ�?�<}�LW1��Y�;n��ߟ�^0����ߍ���nd5D��yß��A���V��>�@W6p��y������!\m'�[�a�~�gX�����_nuY�Ɍp3Ӓp��a?ÿ�`�cVoe`��CQ4�@� 2���`��ĔAY�����7���6���@v퇻�n���e�d��������X���j� ���B?��B���S}���1��a`�W��8]�&��2d�Md`e��0d��HM  ZU���    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:50:59+01:00" xmp:MetadataDate="2022-09-01T10:50:59+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e8ee4c70-236c-6b45-9a1a-ddb69c6b0a62" xmpMM:DocumentID="adobe:docid:photoshop:1338bea2-069a-694d-ba1c-46b590b8c1a2" xmpMM:OriginalDocumentID="xmp.did:17271554-5a82-a247-8125-21b9183e17c2"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:17271554-5a82-a247-8125-21b9183e17c2" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e8ee4c70-236c-6b45-9a1a-ddb69c6b0a62" stEvt:when="2022-09-01T10:50:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Z��  �IDATxڵ��J�@ ����P�E)J���|
��-/�Z<��kjU(z�u)�Է�"b���P463Φ�m�
u!��~��nD$:�o�����o"aah�F�3������>*�׉0 ��V�-	!�C{�Q�	�O78w$�� V��� '"ǭ����S�0��ˣ���  �N�����;��am�ŏ����wP�F�:��7�U3L����8,�P���0��XKЫf1&�k
�Hw���R��a�6�<Bn�l���z~n W�3DmM��*��ɋj���6��s���� 
6��5�������s�m�VT(X��|���j&»_;����#5vVQ���� c�10��NG$�T��%^�D�M�Rj0Ǐs�0?.����߾w����� x1���Dn�VG'{$w�̞;�_���������    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:51:05+01:00" xmp:MetadataDate="2022-09-01T10:51:05+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a599ef1a-fb0b-c24f-850e-e0462e913e77" xmpMM:DocumentID="adobe:docid:photoshop:4e361164-c5be-1b41-83b3-d3d6cff73d0b" xmpMM:OriginalDocumentID="xmp.did:2dc0d662-a807-964d-95b3-d6b8406c1b74"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:2dc0d662-a807-964d-95b3-d6b8406c1b74" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a599ef1a-fb0b-c24f-850e-e0462e913e77" stEvt:when="2022-09-01T10:51:05+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>PN��  �IDATxڭ��K�A ��޹��]��%N�e��"-	C�����V0�-I"�0��RT
�QI�	
$*�b������BT�m���}���W{���s�}x��{_��@���{mmE��'�x��ͦ��5�U��vsٹ{=�Vk��߷<6�g�A[�kWFƝ���9�C��gf������n	l�|l7y��(�T_g3���B!�y�T$	s���^��C1g(#��|������eee�TUV!�=�RPԮPP��1/�����/̘(3�w�R�q�x�#چOVV�,�}&�5P�����7o���T��P�8�+���g���kzv���_(˧��o�h�B>��T����j��Ԭc�}O �M�k4����k��z��C!*Z\Ǽ����Lʆ�ؼ��s���@E���5Pw����059�l(����W��.oq8>k``�3j � ��:0@G���`4 H��;=0����R��"S,kq6}����\�;��\��X�>��;�`2,���5�:7��N��R{�QY&���~�!��%�I��8�_��HVvL���$�6U����{H�M^Zt�T�y`����27����}M	A��Ħntc�X�8�fôM�c #�������ç90[Gl1    IEND�B`� 
BackgroundclWindowNameOpen Workspace (reduced alpha)PngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:01+01:00" xmp:MetadataDate="2022-09-01T11:06:01+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b5b38760-7ca0-0144-9b50-bf916afac675" xmpMM:DocumentID="adobe:docid:photoshop:70e8b403-62b0-304f-b31b-a60a0e122a8f" xmpMM:OriginalDocumentID="xmp.did:e402d701-3891-e647-ba5c-596e1423d132"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e402d701-3891-e647-ba5c-596e1423d132" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b5b38760-7ca0-0144-9b50-bf916afac675" stEvt:when="2022-09-01T11:06:01+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�^�|  jIDATxڭ�[kQ�g��$+*�6�6�IZm�>y!^HQ듖�XA����wP*�[1_4QQD}Q�� U���4��R��I�7g��Ms1���������Y��80��W���F����A�`��������������}�n`,�.�;Sx�l?��<˭�j�]�Y
̾l����W �,��Ɂ$�,E��y9����#���c-,���;C�,>��k�z^7pAJ��)�
;jY.Ơ�ݾ��[^o� �Su�E���lrxp3k�wz���EU_�L%�`@����w�~�ɼ��B̪�	 y�H�T�U�R��o�+ʀ��4`
:�ZV����Z�eE�3H���C�f���nv�/�V�.� ����6{D��(r3.>qc�[�v�.�E�֬�t��|���oc��c7�F7Ht5�:��7W��4���->���S1&%4x�����
����g?�5ɇ��i�m�{�f��++1{f>�-yŮ�)���L2;�����3R�]5��l�i�qS&P�h�,�L*4W��[W<l ǆ|����<�TTRnR��Ϳ5��kD�):�u���ީw�=����x����t%���;�    IEND�B`� 
BackgroundclWindowName"Open saved session (reduced alpha)PngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:57:55+01:00" xmp:ModifyDate="2022-09-01T10:52:51+01:00" xmp:MetadataDate="2022-09-01T10:52:51+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9a883c0a-98f1-6b4c-8769-04ba906f517b" xmpMM:DocumentID="adobe:docid:photoshop:f407ad62-af54-0f44-a94a-c09127aea8ed" xmpMM:OriginalDocumentID="xmp.did:cec3d8d7-80f0-da41-b4a6-0b700ea0fad2"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cec3d8d7-80f0-da41-b4a6-0b700ea0fad2" stEvt:when="2022-06-27T15:57:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9a883c0a-98f1-6b4c-8769-04ba906f517b" stEvt:when="2022-09-01T10:52:51+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��v"  vIDATxڭ�OhA���϶-��H��l�ƨ'�֠��zQ[B=^գ"
T�`�("�^��Z)�7-�[�+bS��i�H����}��$�M��ޛٙ�|�cAD �@�q��f�R꥚,�Ʀm�IR	�Z�����:�T�F��(�M<�������P�	)�\����~e�K=W�ɾcY���)���'�������
!�<#E���_���Hg�����,���1�2�4r�թ�g{�\�(ՄXm�N�.����0��D�`5��P�R�y.�[��M`�28�L�h���9
�}�ec ��}��c>!��P��F���H� ()f� ]� ]&��Y�T�r���� !�� �r���C�V�X��ܤT�s�҈�W<5�p�,��U%����o�}�1E�}�s؏���)
ۢ���D���]��j}�́�O���?R�C/[�bϬ6]�w�M����� ���B] ���2�����̿�����̼6��I�*��ZՖ����	L>ހ_�*l�tg�Zٳr������A�]p�Q��7��lc�����ڿ���ɇM��1uހmI��RX���]����y�����5w���	�:XO�5�ۑ_�M�������|    IEND�B`�  Left� Top�   TPngImageListSessionImageList144HeightWidth	PngImages
BackgroundclWindowNameUnusedPngImage.Data
{   �PNG

   IHDR         o��   sRGB ���   	pHYs  �  ��o�d    IDATx�c���?5 �A��4jШA��A AGѡ�P�    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
b  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:05+01:00" xmp:MetadataDate="2022-09-01T11:08:05+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9e857cef-dc8e-be46-ad20-6937b4c2ebd7" xmpMM:DocumentID="adobe:docid:photoshop:8601866a-4c2c-8d4e-98f2-b3870441e385" xmpMM:OriginalDocumentID="xmp.did:07703220-488b-fc4a-bbd4-c16348e0694e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:07703220-488b-fc4a-bbd4-c16348e0694e" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9e857cef-dc8e-be46-ad20-6937b4c2ebd7" stEvt:when="2022-09-01T11:08:05+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>Z҆  ?IDATx�c���?-#�,�0��?������c��@9���M�����){P,�����P!P������B����P1��?�:��?0�su	�����(t�L���- j �`�B�Y��L{_]�0s�$T�:{�otB3�	�R$�0󺾐aΌ)�4�w����f�?��BG�%T���>�a���4�t����k��Gv=rX��1��2,�7Ղ����[\�Ѽ��$W"��$����9K�A������6�H����Rl�T�7g1,_<Ղ����۝�pz=rQ�ͧ�7g0�\�Ղ����;�b���%"�-��S����kV,A������N�X��D6��T�N��2�_�Ղ�������X��E.������֭B� �����D��������Lbزa�������#
�����@C�C��P�"��ƽm2dؾy=�9���tq���a����wn٠�b###�r}���(Gfj"^ps��`��E(�&�Qn��-;����ENPX���`��|�lܽ���`�֍�Y���G�{wl�D�Z �Q��ܙ~x    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:10+01:00" xmp:MetadataDate="2022-09-01T11:06:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:fd6e66cb-f739-d84c-95b7-eef321ba62df" xmpMM:DocumentID="adobe:docid:photoshop:7f4f77c0-967a-ec4e-b48e-be0adc9f4ead" xmpMM:OriginalDocumentID="xmp.did:0f2d0182-2614-614c-8d72-1d030f1ed156"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:0f2d0182-2614-614c-8d72-1d030f1ed156" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:fd6e66cb-f739-d84c-95b7-eef321ba62df" stEvt:when="2022-09-01T11:06:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�,�>  �IDATx���kQƿ�Wk$��Q�LJD�Y1mƅP""�&�U� 1�\������?ЅQ[�
"�R7)��G ڔ6jZL��dr���i2�W�Bw��93�~���9�aD��<��%@�u`�����(s���wK��I�m��@�Y�i�\aU����s0/Xʓ1��_�<AV��[6�ȠX�w��#8	�wo�P�ˬ
�^	�N����s([��Ȃ�u�y�S�F�@z��'���/5@�u�k����ϼ!.b$�U�� j��MPz� Dfu��1��=XS�O��B���u7�JT��) ư�����۰�����X��Q��_�G��Hb���'��M�r	�b2�z����FL;�|����y %އC�[r� vwc�YU�q���T@�@+~x����f�T�䦱sFҔk��
��
R����.����Z�������X&��}[�H4��M)��n�& �����/��:I��Ñ�K�J�7��W�g��*2Oƈ�����x��J�i@��{�X�F���0�Cax}�źo�P�W/��[~V|}&�{ CN(����hvpCee��>�&!��G�}��r��?�R�W�v��%L�z'����ʝ0    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
/  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:08+01:00" xmp:MetadataDate="2022-09-01T11:02:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8dcc1edf-ea10-fe40-999a-4a132ce4705f" xmpMM:DocumentID="adobe:docid:photoshop:70aad4b4-afab-094d-89a9-98dd4e7b2aa4" xmpMM:OriginalDocumentID="xmp.did:cf0fee2a-b160-df41-88f2-e5159d137eb0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cf0fee2a-b160-df41-88f2-e5159d137eb0" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8dcc1edf-ea10-fe40-999a-4a132ce4705f" stEvt:when="2022-09-01T11:02:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>D��  IDATx�ݔOKA��Yvmڨ�L{i)�=�E��"RJ�ԃ�$Ń�A���~<��` '��{(�#=c�l���f�;���!�]ޝy~����D�~r? ��D]Z�=�
�)m���T�7m�|<�n��|�V?�Z�3�y�ω�w��,�-�B��E���.� �Z�!@xܴ��i?w.��l\�WŴ �����EPcl5\A^]6�y�G@��	�%@QC���d�hOA(��bl���`�Nu��k
�RY8׹%J.C8:�q�Z֫��%G )'�����.��	|��c��LF۝_�.����)�o�B�����։J��� �8|˜s��ۍ��$�~t�{����ڴ[��!�D����!��Q���3��uφ��9| /�p&F �	Qy�0�����r]8��x������h/�oGu�c�S��������Q2nh��a;5����V�4�r��oK���D�DQ���h����(��~����܏���;    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:12+01:00" xmp:MetadataDate="2022-09-01T11:08:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:55521d3a-a212-6140-8b1b-919139565f7f" xmpMM:DocumentID="adobe:docid:photoshop:d1bc48eb-33eb-7942-833d-09818d64bbdd" xmpMM:OriginalDocumentID="xmp.did:7542a10d-6f58-9648-899d-f590c24c5b51"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7542a10d-6f58-9648-899d-f590c24c5b51" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:55521d3a-a212-6140-8b1b-919139565f7f" stEvt:when="2022-09-01T11:08:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>ZO~5   �IDATx�c���?-#�-0<|��60jo�N[TW]���f�����E��[�1���>d�%�a��yĪ���[pˎ,�v�A·��+=?�oH��� �ZhD�xf��=�`>��S�-�D�� "��0v�� �ݚ8ȷ _�[08���HJK�����S�
;Rɥ)���t(�}�Ok #Я �҅    IEND�B`� 
BackgroundclWindowNameWorkspace closed (unused)PngImage.Data
{   �PNG

   IHDR         o��   sRGB ���   	pHYs  �  ��o�d    IDATx�c���?5 �A��4jШA��A AGѡ�P�    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
�	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:09+01:00" xmp:MetadataDate="2022-09-01T11:08:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:012717ec-9b73-d24d-973c-d6eda7591575" xmpMM:DocumentID="adobe:docid:photoshop:78c2b222-f707-d240-b72b-b3501eeca1b2" xmpMM:OriginalDocumentID="xmp.did:6f1b1a15-db5e-db48-a275-cdb0555818e7"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:6f1b1a15-db5e-db48-a275-cdb0555818e7" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:012717ec-9b73-d24d-973c-d6eda7591575" stEvt:when="2022-09-01T11:08:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>g�g�  kIDATxڵ�iHTQ����hPD�Z���!�����Bs)�M�J��,[,E�l��L��P�((Lǥ&[�ZTLˇ�i��K�Y���>w&˔.<�����sν�q���qH;s�p�s��:��mqq��׹�.\�4f����f�lӆ��}Nd�=@�A�`~蚾'vs���������KW!��ѫVC�	�y9YS@��\R��~HE��>��4�	�^0ٌk�i? �g||&���S\{��jw����s��9���M������j-"Z���N����:*b��{zp��:�.�b�)��j�HF���	�A���h���3�͞�q�^;��Oæ�)�TK���'�54<�)�������Ii�r�*n�Ѫ.D��cQ�?<�G��mnh��ށ���P�5w����,��C�HYP�5�6��)D݅�ﰘBF�t3%�<�������|GR�N6i�Iy`�]X��+/M��f�5욘 z��V%�kkp�LHI;@n�tH�����u R���s��K�ںǨ�z�SY, )u?���A�=�F[�=�S���������P�s�|'M�����������$�#�y�1���q5ړ�p9
ߔJ<R��Q53��0}h'�\$�������,`��r�?��Xfa;�D_ѭ�P��@��,�F4�;������d	��H��Z&�l��P9�r���M.ʊo������z1���
[��BHosP!-b[��"*�k1ӱ��X�l���k���V�V��Yy	�ۚ�D_��W�t���f�����
��?�������������_p��nX3x@q��"���¬I\]-�Аܠj�_��_�;ҁ,��ྫྷ�鯀��~}MacV    IEND�B`� 
BackgroundclWindowName Open new session closed (unused)PngImage.Data
{   �PNG

   IHDR         o��   sRGB ���   	pHYs  �  ��o�d    IDATx�c���?5 �A��4jШA��A AGѡ�P�    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:02+01:00" xmp:MetadataDate="2022-09-01T11:08:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6e1d4c2a-ed3e-ac47-8ba9-3b3e9df2366b" xmpMM:DocumentID="adobe:docid:photoshop:d6ccbe45-8196-414c-a64f-e8def589a2d1" xmpMM:OriginalDocumentID="xmp.did:3b1b3a48-6313-ba43-a818-89582e3482bf"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:3b1b3a48-6313-ba43-a818-89582e3482bf" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6e1d4c2a-ed3e-ac47-8ba9-3b3e9df2366b" stEvt:when="2022-09-01T11:08:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>g3�x  �IDATxڽ��/Bq��\sc���lLkk��ղ��(�RJ$*E�P1�MI&6����q�<��)-?~��9�����s�="�_�߀���؂<|�ʭ�����n��/��򢿕 ��G�L�Z��C8�����٤c��C���D�o �@��@tm���9�[ML �B�H�����[� 2y?lonP�1��)��	 �)`w+J�c
�.@,���N��q'z�N&@�X
�{q
�����q1D�H�R�`�a��fEbH�S@g�`0�at{ }rD�ބ���K �L*A��a�>�|���A���c!�C>`����׃�.Β���r��J&秺�\!Y�/3�fpW��Ñ�q����}+"�q(�����l����#Y���/>�:�_�F�@{��"����:������*������
!Qu���4|    IEND�B`�  LeftTop�   TPngImageListSessionImageList192Height Width 	PngImages
BackgroundclWindowNameUnusedPngImage.Data
v   �PNG

   IHDR           ��   	pHYs  �  ��o�d   (IDATx���1  0�_�P�A�h�Υ�@ �/��_���    IEND�B`� 
BackgroundclWindowNameSitePngImage.Data
	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:06+01:00" xmp:MetadataDate="2022-09-01T11:08:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c5c046de-b655-cb49-9c64-c7c15b903579" xmpMM:DocumentID="adobe:docid:photoshop:ed01a016-66da-ee49-94f9-5358d678a6ce" xmpMM:OriginalDocumentID="xmp.did:60762e20-588b-4c4b-a207-be67be5ef6f9"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:60762e20-588b-4c4b-a207-be67be5ef6f9" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c5c046de-b655-cb49-9c64-c7c15b903579" stEvt:when="2022-09-01T11:08:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>.,��  �IDATx��mOA��>�!���і�BӠ�&$j H����T	)`����-�"����A?�`�[_?7�^w���`���4��߽����tG@D��G�g B��Ҷ�Je�u���O5��hL;.��\��Qm��L<R>:����f������"�y� �͇�s��|X5J2p�<�^��(6��!^� ��W��9�k������XՁ��{�S��(�˹�O�Bխ��x��,�������ކ)��ls�&�p��c��X��� S3s��ݤnՉ�ja��ra��3�}���� ����z�;�\������N7�}��r�L>��-k��]Soq:3��cR	���X�����帡��3�u�w�� �\� ��),Zn7��M�u�e	VSq
0�`�r���膅�]3�����I
��M* w�դ�������L�q����s��_���͵4p?��N����h�7t��E�떟Ȭ�R ����\���X7w��+�n|� �n/-��:N+a�g>Q�1������W�6\Ƈ��_�����w�7q�^�����.�k��
02�B�l�)�L��_l)ƴ���V�<G�v�� �����Z���Um��� G����Sv>;V�9J��-JA0]JG��n-�hxȴu�V �xJ`�����vȂ�u�]ik#���.C��0�\@g��%��b�<�e=�� g!?*o�1�    IEND�B`� 
BackgroundclWindowName,Opened bookmark folder-stored session folderPngImage.Data
e	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:10+01:00" xmp:MetadataDate="2022-09-01T11:06:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6123b322-6c8d-8647-8f82-86944185aaea" xmpMM:DocumentID="adobe:docid:photoshop:49750230-1405-654a-b5b3-f7b1a60aa2fc" xmpMM:OriginalDocumentID="xmp.did:5a3be35d-af8f-444f-b58f-3c89f571b4af"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5a3be35d-af8f-444f-b58f-3c89f571b4af" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6123b322-6c8d-8647-8f82-86944185aaea" stEvt:when="2022-09-01T11:06:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>x���  BIDATx��KLQ���k�-��}h��(�� A��F��L�ׂ�;��r�J�#nLt�EY�R�1�B�P���vǙi;L;3ehH�L��̝����AD(d#��� ���ҏ@�� �pW�����E f��j�g��Ku����s�!�����?f
 �(�H'�O�D�� ßnX�.�@�Q=b�����2��5j�4VZr(HT�R�+���PT�@Uª[<<��"@�2�b��h��(�ʛ�������a�@�����ъkX ��ER�.,��0-�Ė@$��]���Vh� �/dZ).�B�;ll�_,� ���&?������jPE@�'�F\��~s��"���$ �oG_�Z����%�+M�Y�(D8FʆW)�g1QG��	� �gI�����F��ڗ���@�JQ%�u�xr<�Č��Cz
~?M�F�P����W�H��^�U��!S�{���I҄3&��~�le��ʒ�J6��q�,�O����n�?6@sϥ�"�N�5��d	3��iOq���0�ȍ1��հ��X����!��?e�{2v��C7�狡һ�;�5ͣQsz��" 1d���� ��qra���-E:�Nk���i�E ��������N��R��yV�D�4��-8��@�^[5x|���
L���N�6�2�Eg�XW�)/�k��-�;�����[U��q�C�{�JI2<��98N�( >߭A��6(-�����l�Z/,���?-��( ��o��m��|����9Dr�s��7a![��FH��ɔ��    IEND�B`� 
BackgroundclWindowName,Closed bookmark folder-stored session folderPngImage.Data
l  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:08+01:00" xmp:MetadataDate="2022-09-01T11:02:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e7bbcac2-09c2-9741-bba9-a721dd2243cb" xmpMM:DocumentID="adobe:docid:photoshop:d839a3d1-87ad-2f49-98b3-f353c535cb1b" xmpMM:OriginalDocumentID="xmp.did:733049d7-dcc9-644f-864b-ee70f7c2ee15"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:733049d7-dcc9-644f-864b-ee70f7c2ee15" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e7bbcac2-09c2-9741-bba9-a721dd2243cb" stEvt:when="2022-09-01T11:02:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  IIDATx�c���?�@�Q�:`P8��^�	��r�302aU������v�絔X�ͳ`��#���(0�:b-��{�4Q� �w?����~�b@@.`d���?#�TV�g9��[��Y:�����T�3��p��I{:#V��,��LL��b��?��3ÿ?@s���06���ȁ���W��Io	v����W��G{Z�������5�r�e��B�cd���l{	����/k^�Є�d������� |����h����H���b�r�`�Y��Q����8�,��a���(V�{x`��#(��o��EOt�e�:?�� �t�f9������<0J��j�9
��X]��q�a�
W�b�A���bQ�yS����w�~$�Fl���G�!���ð #(Iu���Q��_<Y��F���:�Dd+\�B+���xh�,ˉsv�	;@Ӄ���?�:< � ��v=q�?�T��<�ܢ�W���_��#�R���>8�@zP&���19 �&���raO�:` ��;  �� �h��s    IEND�B`� 
BackgroundclWindowName	WorkspacePngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:12+01:00" xmp:MetadataDate="2022-09-01T11:08:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:4a716ae3-7016-ca4c-ba15-43bc1da6a3d5" xmpMM:DocumentID="adobe:docid:photoshop:fff55d68-7635-d446-a82e-c7d2e2ca642c" xmpMM:OriginalDocumentID="xmp.did:690ce4db-4039-2c47-a9fa-4711a18024d7"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:690ce4db-4039-2c47-a9fa-4711a18024d7" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:4a716ae3-7016-ca4c-ba15-43bc1da6a3d5" stEvt:when="2022-09-01T11:08:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>ѓlU   �IDATx�c���?�@�Q�`t�✕2#�z{o�.9�A���ڀ8������.�n��B0}ּ���^X��p���@��r �u�6�̴�A�  ��a��v�v�-;0�v���p H1:��'E����� �)"`zkΛ�ထ�!����ထ�K/���z��#/
v�� �nM��##
$�����O��"� �IF7��v(�;` �� }|a���U�    IEND�B`� 
BackgroundclWindowNameWorkspace closed (unused)PngImage.Data
v   �PNG

   IHDR           ��   	pHYs  �  ��o�d   (IDATx���1  0�_�P�A�h�Υ�@ �/��_���    IEND�B`� 
BackgroundclWindowNameOpen new sessionPngImage.Data
�
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:09+01:00" xmp:MetadataDate="2022-09-01T11:08:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:49f9d9a8-3235-5248-9683-b9d661b9c32a" xmpMM:DocumentID="adobe:docid:photoshop:e5817a1c-7f65-4041-9b6b-87c00693b026" xmpMM:OriginalDocumentID="xmp.did:bfeaec89-eee2-424a-bad6-3fb92e9e84f0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:bfeaec89-eee2-424a-bad6-3fb92e9e84f0" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:49f9d9a8-3235-5248-9683-b9d661b9c32a" stEvt:when="2022-09-01T11:08:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>C;/.  �IDATx��{LTGƿ} ��Z��)��	P5��1iL[��(%����#Ii$�P,!�Z-%Hy����(����6-�mڦTK*���X�u��ew���J0���lf�ٙߜs��B�XV����{�z^�/��I�;�h��Y�WT}�a�w�bX7�0�55)��c
��dl;�a��a��sۖ�I����� *������#���q��lљ�@����>0��&;��.j������3�x�#�DE@�^@euJ���q<��k8WR(� ��ipga,-�݈�1Û��SD�ؽe#�n~�h���?�v@�Vݫ�5��p�l�WPD�"��7�o���h5�37wF�U�^k!�ޡ�pq��Ԩklf��!��"�H�0L����B �6-��f�ð�����>@X�?\]]������K�9��n�F����E������ޠ�p*��4��3'm^���_<RȜ;\777Ӧ��e� K�ޠ�/���B1���B- 'O��(���� �1�
>�M���������oS�-���Aϭ[�Q���W�MNN�� �~�GZ�yQ�>J����L#X�@\l��ds[���_�����K_�A���i�c���n���I{���"������[s�@�7ߢt�El�AU�E ;�i����w��&��z�V�#v_����E����;g1�+ŵ��4@V�I"���]�����x�K��];�A8�f�;w���c̊�E�TBv�.�o�PSUA���%��v���±�[�1$n[�M���OP�ԐͿ�7���k�c��p��7:��w7Q{�����a��uG9���@�~����DÔ��,��{k��eLNN���T^<Od��&7����ǧf��i�t�B�Fun6�E� Y=	oW�{Zq��
��q�����J��F�uc�u�==`�Һ -��)������X�m�w��������HM�$]��e-h�y�zzZ��K�"�N��e��%ئ[N�9J�OLټ�[^���z�Xj:�$П\'s�U�������b��Hi��)iĚ�l�]N��>����~G[�ѱT���߅�d�r�,�����)k�><z\��1l�Nʝ�3�9��.Y3�(}�g��Ğ�����o�e\�t�.@���g���Am��Ą�yT?r_����lY1����0G�S �U��_�ؓ-i�    IEND�B`� 
BackgroundclWindowName Open new session closed (unused)PngImage.Data
v   �PNG

   IHDR           ��   	pHYs  �  ��o�d   (IDATx���1  0�_�P�A�h�Υ�@ �/��_���    IEND�B`� 
BackgroundclWindowNameSite color maskPngImage.Data
E  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:03+01:00" xmp:MetadataDate="2022-09-01T11:08:03+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9422131d-8f21-b146-8f19-c722622a2620" xmpMM:DocumentID="adobe:docid:photoshop:4abac5af-6043-9844-a8c4-fc3cbee843fe" xmpMM:OriginalDocumentID="xmp.did:bf469140-3c07-e840-8257-dcbfe1d6bcf4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:bf469140-3c07-e840-8257-dcbfe1d6bcf4" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9422131d-8f21-b146-8f19-c722622a2620" stEvt:when="2022-09-01T11:08:03+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>x���  "IDATx���Qo�P �ӟ`��|�u�m�͉��c�b�6�v@Wk�!��nBpnFs�����8�1�gb$8�|�Mڜs���M_��p���o �l�ݍ�;�;��;�~�s����k�s��X.�29� �[/��@>���Le1"�2V֠��P�am��4���B1���3��g<���]����RT`x�h��o) ��(K&�ť ��h	Yd�x�P�*R�����Ę �TJ6(Z��%���S���1�Rf���Ze�$E���p��v�e
��*�	�	�Μvk
%]c��]�O;U
�De4�8���<�wk ���z�`������
�#1L�֙ &n�B�����)�	�ƭ8h�Q@�������9�f��a�mӀ�j�Z��r�b�ؙ>hP�r��ӽ��p$`���}���k�ʏ���><������M�띵���[��)�8n�X�K{��oq�M����+>��� �#rී���.���|����n�W�aǙ��&F����k\ �AK�ϻ��    IEND�B`�  Left�Top�   TPngImageListActionImageList144HeightWidth	PngImages
BackgroundclWindowNameLogin (reduced alpha)PngImage.Data
(	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:07+01:00" xmp:MetadataDate="2022-09-01T11:06:07+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:158c467f-8bd5-b747-86ba-c44ca85581eb" xmpMM:DocumentID="adobe:docid:photoshop:1f376027-3424-4e4e-85ee-c980b18d4d7f" xmpMM:OriginalDocumentID="xmp.did:9b2376a2-de62-f446-bd73-41c935f71535"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:9b2376a2-de62-f446-bd73-41c935f71535" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:158c467f-8bd5-b747-86ba-c44ca85581eb" stEvt:when="2022-09-01T11:06:07+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  IDATxڵ��OA���H�RZ@��Q(��h�p����'߁�����P�/�Ah�?�%�*L��4�-]�E�Y�*	�i�ݙ��~��M)�ap��� k���B�m0�A��.ż|_�r�Jڴ�.�Q����τ�N2�o��p�ڗ)h�1	��!'1�X0ؕ�=���H�?�`j�w�ZNE(fA��<o���" #2 �BFp#�J��1��?��o����&x}Kp����Q9p�OL��6��U.�}�E�i���A�*��Ɂ~"׶S�(�1��)����ӽ'�r��e��+.	�Γ\=Q��:�����.�C;���9vȀ�5곝 v�ʸ8�W|�fі�"����m��b���F��z������� ��XU"$ɀIS�04�-4ù�F���u����y�d@r��O��t���f�D���|�qf����<�?`Fr��pȫ� +[OVA��'E�b2Eߚ���)j�R>���$���u���k��&�`�?^�,4�41��\�+�6<�(�QS�����v�{���f'�,P;$D�6%rh�Z�od�J��롋J����m���p {��"���F��U�A��|�P��R O j`}Zd��M�c\O��{UV�B\��1l��^BM��ȁ,��ez�wO?GX�r����^���P�7fe��,A���'��޼�/R��2���S)ע}�l?���y�\�W��U�EQ�u`�>�P�W�v�=��������@R    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
�	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:13+01:00" xmp:MetadataDate="2022-09-01T10:57:13+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b7ddeec5-6134-f84c-839c-c49e418fe837" xmpMM:DocumentID="adobe:docid:photoshop:a9fd7f0d-1f94-9d41-a78d-ba83d2cf4320" xmpMM:OriginalDocumentID="xmp.did:37df698e-d87f-e64e-aa08-743c8c3e27f2"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:37df698e-d87f-e64e-aa08-743c8c3e27f2" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b7ddeec5-6134-f84c-839c-c49e418fe837" stEvt:when="2022-09-01T10:57:13+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�'j�  {IDATxڝ�ilLQ��w�,-��Q�W�D��"�D�R�'�D�H+��(*�V�-Em	k,��K���� ��%Z[M�̴��-�{oj̛ż��͹��{���s��=m��� �A!�]�6����v�s-�]�%�V�������.+?s4`�w��Eh��K+���u��p:y] �;�n;�PX��V��S�/��}HH�u2�f��fګ�� ��;h���>q|#��1.�5�`gGN�QL�;�����VO�P6��8����<n���66���?��r�
�ԅ�,<@����� ����6S��/?��'�6��ѤTY�J�c@��A��t\i����M{}<2��j���`Wr�V0�h���	��֎�/g��C&XO|s�x���� �T"�T���6,H�A|,�N�8��<���˄��!��Q�p"J^�>1z^�7�SB#���aQ[7�&8�&���R�.�Ɣ�p? ND���c*�0�(�(�`���:��u�ŵ#U jds��Q�H(�߆J�J�$F�t��(���-V<m�K�c�Ҭ��$�"R�Sz7�y�S�m`�/��"���7�Z�`G=��;{�T��D��.Xs1:��眕��i����N8���N|����GD�>VIā���Ry��F�|Z��-�]�t>b����-���EA�&�r�e/f�A�J|�X��Q �k�OD�/�F�ݰ�֎�JpO�	OdJ�x��,�V8=f��ʯ�E�^�����ls)���Q�:�>e�� Uܼ�b�z�`�y��t3t⾽��Ɖ���z�?닊�5��V���"��B�s�9 ������FubD@�����?�p"�҂6�W�U7��x8�`ʌY4��@ii�p�
�B�    IEND�B`� 
BackgroundclWindowNameRename 2PngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:15+01:00" xmp:MetadataDate="2022-09-01T11:08:15+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d36b3ed2-f4e5-fc41-87ad-ccc21c20dbb5" xmpMM:DocumentID="adobe:docid:photoshop:c1b2245c-e1d7-7c4b-bf8e-25710f5695ac" xmpMM:OriginalDocumentID="xmp.did:318a5968-8b6b-e040-a2ba-0cfc71cc5cd3"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:318a5968-8b6b-e040-a2ba-0cfc71cc5cd3" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d36b3ed2-f4e5-fc41-87ad-ccc21c20dbb5" stEvt:when="2022-09-01T11:08:15+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>B���  vIDATxڵ�YhQ��$��6�"�P*���F��U|�D4R�}�SQۀX|��)�!R�"(��}���E�ZѪ)UĸŚ��,��q2�C�1m���e���ߙs�P�  EQ��"m�=(��S�h�껉))[-��6�FB�l<�ac	��cuA�Stk�>KO=���Y��%�A]5��y�h2;�rZ��!�&�"�A�b@z�Q�g��fK��{�3�<�_wy£�Ș�>��;���|��ߢ)Cr[[Z�q� 4����7bq��cw��˜+|،����3+�,�� ���cΣ�G���Ȅ��8!b-����b ��a�ѸX�N��b�]��\�?��As|��1��s�@���ݶ8� <��C������fzkx�Ooр�Ȧ
�M��1g�*U/�%�pk>�8�h��Z�K�r@,0H�?���{�R2@|(�x��ֈ ��T徼v1s> �R�s��*�g�����Rh��ZO^@��of>��*�+�d�f�	t�C eu ѷ�����\����];Z���!�?^������,�^�� ��a1x�>0��_0��!����N�,1-*����y Uӳ��S?������J    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
A  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:51+01:00" xmp:MetadataDate="2022-09-01T10:51+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:cab01aa4-2548-5d49-8eab-9e84e5623de5" xmpMM:DocumentID="adobe:docid:photoshop:cb0114e1-8033-a04d-9949-32bd9e4d032d" xmpMM:OriginalDocumentID="xmp.did:c818f13d-6239-1d4a-a6e8-292abdef8f96"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c818f13d-6239-1d4a-a6e8-292abdef8f96" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:cab01aa4-2548-5d49-8eab-9e84e5623de5" stEvt:when="2022-09-01T10:51+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  'IDATxڽ�OO�@����(���1�$ {�1	1&`��J4�(G��p���	�{���~��B4$��z��vw��x3m���5��ݦ�����f�F��	d*���[��ߜ~{╅7kJ�;�w?��&'�P�[|k����n(�H�4k.�T��J����)���s넸��|�R��Ix�O���L��}{Uw����_��\IN��bq��������g����%C%�7ޟz�$#Y��#'��Ι��E��y��H^�v	��srz~f W�	t;y>Šˑ�P�/����du�U��h�;^J�ě{8ѫW���LF��p�w���7᱓�ɀ�!p���&L	w;$K&9�H6�G����k�%�kW�ǔ$W��h�M�ѣj\�QN��zA�%�?ъ���yy��	h��v��s#*���R��J1��7̲b�x��bq�ҋ����:m��'�Ӄ�,A'�2PО������>V���_���[�Ҙ����}ux��^7��-�Tn.Ll*�,O��Re��~��~/�e���\p���C�h    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
l	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:51:06+01:00" xmp:MetadataDate="2022-09-01T10:51:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0ffffdea-2e6f-c449-871f-3061b89845c8" xmpMM:DocumentID="adobe:docid:photoshop:71b5c369-cceb-834b-a39f-00072bf3ba76" xmpMM:OriginalDocumentID="xmp.did:a2732e9a-438e-8a43-a90d-b7a9c528e5fb"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:a2732e9a-438e-8a43-a90d-b7a9c528e5fb" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0ffffdea-2e6f-c449-871f-3061b89845c8" stEvt:when="2022-09-01T10:51:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�*�  IIDATxڵ��oQǿ3�AV��Z����Dm[Ѩ[� RE�{[�l�ċ�DB�4A4DD�K	qIфͪ�e��Jw۝��9�ݎ��M[��L��w�|?�˙���8��8z��z�c!94}gu�+�=������>Xm�1�ݞ�m���S����S���ue��s�?z�&�v8Z�������y�b�=MM��WNW�bk@l4�;�׽2�о���q�dJMo��Ƴx),5x~ú5HJQ�2I�D����C<g�� ·�R�yLׯ�+u|F�k��Y��e�E�` ϖ�$C��],��`�0�A4=y&y;:�F2�m����۝��X�x)233cb�2E ����>�C!����j�s� ?<��0$㓏C�s��/DFFzĸ7�	����0�������Q{�~ɚ����3`̚	
��D? �p�L��6kV�T��(�t��5���(����B|�����ؐ�U}+W�d�oARP1g��_Z�s1on�Z�����hmk/�uT�Q�z٦�`���$1��z��l] �5*-�gph��b����x<p:��U[�T��V��D�(bHZs���Ts	�2���z�7�9).��v�t --_�v���ܜ�L�RI�+���}2taRj3.]#"(�K�L4�fU�TW��
�#?���(ƿ��fY�Q��_�)��2P��4�ӄ �䵚�h���Q\��ս�P�Jo�+AbM1��4#1 oEL��i6���/�옾�B	5���r�	p3�%wa4Rq�6u@����dLɀ�4�߲�4MS����<.�av���?a0�S�=�ֳK���~���6=�s    IEND�B`� 
BackgroundclWindowNameOpen Workspace (reduced alpha)PngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:01+01:00" xmp:MetadataDate="2022-09-01T11:06:01+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:2a0248e1-0d38-f649-8980-e97715a22ed3" xmpMM:DocumentID="adobe:docid:photoshop:4884fb40-fb21-3141-9aae-cd073f5d17d3" xmpMM:OriginalDocumentID="xmp.did:8bcd2802-ca77-c941-9b0b-7a7a4d752f88"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8bcd2802-ca77-c941-9b0b-7a7a4d752f88" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:2a0248e1-0d38-f649-8980-e97715a22ed3" stEvt:when="2022-09-01T11:06:01+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>X�m�  �IDATxڵ�MhA����TZbm�X��hŨm1m��VJCQ� �

��9	���xS��b<*z��~U(����j#����b>7�>gw��&٤����7;�~���w�c02��a	�~���b ��K�j)�~��\��E�xq�ı�'�]�ƭ; ��z��pT�~���c;+Ԓ�$HY���䅲���~���k	���,�D >�~�
p�Yԃ;���� �X A����_� ��)���5@�j+�v]b?��$(⛈���jK"(�3��r�*��+5m��|6�Ae�%{CR���b~% ����3H�@�%p���z4lu�f�&9bj2_(/ ]�?��&�T ���1`ԛ��y���g/���U�q6��h��;(��j1�'��qg��Ť�1�Hv�������BUѼG��dEX����y�Ԁų���F4u?P����ԣNh�Eh�N��%e���0{L���S �49W{�T�k�*#�|F�!%��J�������t�ܚ
�h�)[M* �82a�텤 ��S X�掃�X��5`l����)>
�������-����X0;��#y����� >�o�z�u�D��u�P���^�w�Y����L�kа��OJ�+#X ��ͻ����Hd S�>�7�'���N�7�5�a�;3&�Ӗ����<-s�    IEND�B`� 
BackgroundclWindowName"Open saved session (reduced alpha)PngImage.Data
7	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:57:55+01:00" xmp:ModifyDate="2022-09-01T10:52:52+01:00" xmp:MetadataDate="2022-09-01T10:52:52+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:1c12d99d-a821-6647-b7d2-2bc3ec89f991" xmpMM:DocumentID="adobe:docid:photoshop:0aa16207-d95d-a843-a727-d6870317f6d0" xmpMM:OriginalDocumentID="xmp.did:359403e5-bb6c-554b-9564-ddf6fad1bf12"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:359403e5-bb6c-554b-9564-ddf6fad1bf12" stEvt:when="2022-06-27T15:57:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:1c12d99d-a821-6647-b7d2-2bc3ec89f991" stEvt:when="2022-09-01T10:52:52+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��B  IDATxڵ��KQ���k-�i
�X���h�� ���,����?�܈�$�
�R$*B����TZAۋ!�C�d���/tם��{�;3���ٵ5h�r�;��9��3�r��A:�����L[>rDY���hc��9�ͭ
N��h��j@�m���X�%/��uò M�o��*�ND���q ¾�;��i����ڸ��$R续���V���L� ņ	`륷?ϵ� 9u����3xo���wSD���Dq�wz&r��p��k�~���=a {|�Z}<��"�����@,%��=����#5 �7�	:8����*hZ7��/� x�^ >W�&�L+!��6�ӝY��{	h��&�=����Q�o�~���m06��ˏC�-O� � �0��&�0��0@�)P�����!;ST1��*�E{�6�h$ɥ ��|�g�O~*�σ�l�/dmh���K�Y
`�	�"��'�j<�\��A�?`�k�A�n�C�>�q�A�d���C�\ƁKG�ڜ,teT6(��<�/@._y�v}�(�M�s�b���ץ &{�qd�[*�-+g��H��dёHؑ��*��;�
��ī I)&���& �.���=��h�N��7A��H�RL���@a������1��
䬹`/q&�<6�b��T�6���8�-��r��4�>�D�2"\�w�Q��-�5�v��Q�X`�h�@�v?,��� #��6z��X�NH��'N��X���%i]��߀?�̷Ƴ���    IEND�B`�  LeftTop�   TPngImageListActionImageList192Height Width 	PngImages
BackgroundclWindowNameLogin (reduced alpha)PngImage.Data
1	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:07+01:00" xmp:MetadataDate="2022-09-01T11:06:07+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:eca146db-ddec-7549-98c6-7d2cc83c44af" xmpMM:DocumentID="adobe:docid:photoshop:8cc12f2c-50b2-314d-86c1-47e7ccea188a" xmpMM:OriginalDocumentID="xmp.did:e46918be-2d69-a347-b630-d628ef05a718"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e46918be-2d69-a347-b630-d628ef05a718" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:eca146db-ddec-7549-98c6-7d2cc83c44af" stEvt:when="2022-09-01T11:06:07+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��6  IDATx�͗�oA�g�hbL�-�_|2�w/T��d��j�O&jS�S�Ǔ-WK�I�j�j��V�>e����.���1��b�f���}���AA+�� ���1�h�B��9�4���
�3.�j ���,�wV�ڑ"����X��I�R���C�_��knx�o�9�v@����:���� z;jh)�� e*���׀�3
8���
* �#��W	�"`s��D��6\q~����,�>���j�cnK������'c�W� t��nfPH��xFƲz����C �듌�<��Qh�F�[{��	��t O݂P?�B@��* ��I>F�P�� �Oxc`CV�,
1X񃢤m[� OT
0��Ai�*EVcje$3F5"G� g��[@�!b�:K�E�#�EV�Ǜ��1�H��pP���1�&jL�t R[��	�~�4�3V�+ #	�@��q@$�5 g=�Bԓ3��C��~Q;#�R��d�� (k]8�@m��f ��Q������.�Ǝ�ؙA����ʳ ���Ԡx!%\X�Z�˺�uc��(�#�X {E�D4�])8���ڢ'�}�'@�h �|�dI�
գ���Q>3 ��"�s����<� ��� ]�50���?$Pz�%�qa��Ggz���&�mi
B>�-n/�����[��`�Z�_i��#Ŵ �l��b_:�t1ٸ��tn����������M�_�]LjW3�t5�k|5㤫Y�r5kUi9�_
�u�1��    IEND�B`� 
BackgroundclWindowNameOpen current session in PuTTYPngImage.Data
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:14+01:00" xmp:MetadataDate="2022-09-01T10:57:14+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5a533d10-ab3e-d942-9287-314091b55f5d" xmpMM:DocumentID="adobe:docid:photoshop:6014b440-d073-5f41-81ab-c04801887a2a" xmpMM:OriginalDocumentID="xmp.did:0a34ae79-7d96-5b45-9032-45160dbeebda"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:0a34ae79-7d96-5b45-9032-45160dbeebda" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5a533d10-ab3e-d942-9287-314091b55f5d" stEvt:when="2022-09-01T10:57:14+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�2�  �IDATxڵWkLU�fv�݅V(m��4XJb���?|��R�h[5E�4�4�RQZ*}Y�����@4Q۴Fc��@�h���ey/�;��ݧ��,��t�7g�����{ι��@���x�_��8:�4D�EH��m�g$�6��@}�Qr��4�O(/��@-�.��O��PE���9���r�`�s����3�Ϩ#P[w�\Hɔ���2<�Ha��(�ߏ$��{N�#PS{���e����JM��\)֓>d�q��S�AFO�:U5�Ki/(�j=ߋ}�X�T�uz[fOa�������s=����:@ZS���I�*��D�"A��2�A��R:7b�'�(��"m�/�&"��l�	98�������»ŸfOZ�����#PZ���o��D'�P�B��g��j 
"��ّ9�x�U�����c���V�+)�#�`?W����0D��/,(�NM��%�N��?��S�jTG�����IJD-_�ez:C��q�;�1���'1�,�y�A��#�|���u�F�Z�0��08���uȵ��^��I��C#PQ���U����tլ����vzr{F���Lb@����t=��
���ׁ���a�� �$���Y|��ڤ��ɮ���!L_[f1²��A��� �ޓk70�#��f����V���uA�E��yh"m�G��B¢hw"�����[tt�I �Ӯ(�mD�]� �������K+���hǐ�ɠ[�������Ѕei�'�b�xX&9��f�k�m��j�YHX��P�)�h:4��F�fs`l6��w`e���	�',J�;Is�Q������a�ʡ�_=��1e���:�/&,���KS��t��,�43.p^��G���/�[��f��E1�ߣl7��@�uW�7�κ��	��I������f��m�}ڒ����νsWY�a8}=%:BWX|P8�9�J�Uo LC|/S��k4^�-���;q����	8��#啠U�-�R�Q�6�yVp��d<^�)�ٶ�%,__8:����Ig��`�dō��X����y�e�	��큃g}����U��
�HW��y��oF^Dq�����ww�a +@X�im	�@n�{D֯���"�m��dt�Ʊh�����(,W�U�۹�7%"=,#0����Q��X9-j�}��ea1�:/�%�L`���h"�"�"'�-U��	��u��ژ���G������}!캯�2�.H@IX�\��O�x�%L    IEND�B`� 
BackgroundclWindowNameRename 2PngImage.Data
d	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08:15+01:00" xmp:MetadataDate="2022-09-01T11:08:15+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d7add81c-694b-7f4e-a510-1f6e78dcdbc4" xmpMM:DocumentID="adobe:docid:photoshop:a3b56b8c-50dd-b64e-a16d-8057b168c3cd" xmpMM:OriginalDocumentID="xmp.did:075f022d-11c2-1d4c-86c5-e6a33aaa9782"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:075f022d-11c2-1d4c-86c5-e6a33aaa9782" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d7add81c-694b-7f4e-a510-1f6e78dcdbc4" stEvt:when="2022-09-01T11:08:15+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>W��<  AIDATx�Ŗ[HQ���]g5�55�+�փw�
ɲ��$#l�!��J+I*�*�J=%X�C���J�$I׊R��l��Ι9ӌ�����e�33g��}��B �cY\%F�Ym�"��Ϗ�����MU�dkc��� ��<Bv�<���T��e+;9�MCv ��H|���ϔ]������˛�Gu��p0�K�ˉ��\V��FS��d2�X�\�x8�E�FX���	fY�߯��T�A��B�X�	��Z"�W[���7���wԞ�K����=?�*LV6�d6;<��`Gq���~�޼BC/�Ƙ�̂�#^;[���,E�7��*�wd��'�����⠊�M���r�&�hώ��3��
O}��zU��
`m�ḳu����c$.����̔��#��๻�\;GA�C��w�/�g���5���^�ٰ�KpB��0�)�e�7�vOn<$}�Rj���l�>	���l�m8D�5��L�~mu5`���A�N��Ql���o.�	�8����C�\��Z��f�g�O\���?2�u��wd.Wa^l<��D�?�H�(��=�z�0פ��g�\K/����'xT��{K�	�f�4���LM*=�����E�T�É�=����`$�#!@��$x H�9- t��.�&u]Z&���]�
R�KA��2J��+d�CW}�g�� zk# ��_�G{�k �f�]CBx�!��P+��c�W�5hzo���~(*;�q�^��8��,vUUU���ܻ
�����@���Q`�m�Ϙ��S��	����`���y�    IEND�B`� 
BackgroundclWindowNameDelete filePngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:51:01+01:00" xmp:MetadataDate="2022-09-01T10:51:01+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:41d20d2f-3c6e-aa43-aefa-8e9d8b8a72b4" xmpMM:DocumentID="adobe:docid:photoshop:1440d40a-71fb-8b4c-b619-25e390ff0d7a" xmpMM:OriginalDocumentID="xmp.did:df096d51-cb03-884d-b8f7-36e4beedca68"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:df096d51-cb03-884d-b8f7-36e4beedca68" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:41d20d2f-3c6e-aa43-aefa-8e9d8b8a72b4" stEvt:when="2022-09-01T10:51:01+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>\&�3  lIDATx���j1�o��"-v׵���σ�EzQ���P�>B��w(�"TA�>���h�ֶ �X��I2��vg���Jo���0��MNr
 �2�p(�����=!�l���A@~�ԘY�V����</��Xǒz*����u�h��
,�\�R%�7�v*I���|9@�?����oN#��ƛr]8�t�գ}8�3T��w�
�6�(��%Q���(.�����	�����x���Ӻ"-�2�#�?|G�H,gK�����mF�
 IGi�>��W���/n1 ��;�91��H����/-�%�P�R���� ����+	诜�a8p$���xe-1[�pP��F�0�(��M�p�?�:m���Ep;"�y�����C���f�C���M�\8�\��I� ��U��<��|���v�mN��]�
�}��/'��ܖͩ�'ܳ�y]�Ix	��۲�l�ќ6��'��Qܾ��7&����m���Ɤ���+A���ܐ�%rv���S���:c:p�,~�4�H�}f\5`�p[�=��pPŹ�?\��}(U!ؙ��Q
w%Hr2V�G�g��I�==*���Px*�xHX�
n"�#p�J�������Y    IEND�B`� 
BackgroundclWindowNameCreate directoryPngImage.Data
�
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T14:09:55+01:00" xmp:ModifyDate="2022-09-01T10:51:06+01:00" xmp:MetadataDate="2022-09-01T10:51:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d88edd5d-346d-d74a-bc89-2fcadaad2ee8" xmpMM:DocumentID="adobe:docid:photoshop:29631f50-33b9-0a4a-bad3-40c6be495783" xmpMM:OriginalDocumentID="xmp.did:e7313573-7b2e-7f46-8b80-c48a2837d230"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e7313573-7b2e-7f46-8b80-c48a2837d230" stEvt:when="2022-06-27T14:09:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d88edd5d-346d-d74a-bc89-2fcadaad2ee8" stEvt:when="2022-09-01T10:51:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�B��  rIDATx�ŖmL[Uǟ{��Q',i� ��9&Dcbt�l��+��2$V��Lf��?���3��dD35�,1s�aX�n��X
�2֒JKo��r<���޾\n����s������<Ϲ�@A������|�^1� _�l~3�<�����罢"s��9A��k;���W����,,*�66�n��b�׮�>��K�+�s�w�Z��۳��������!&(���Y��3���T�-8l�����7�:��+�m�
���c������\�,��=Rh�*��,Pp��!�+
/������ �`����1
��O ���눰��O?Q���nݬ�h4�ŕT��T*q"�# ��� 
ò@Q8�0zs��0�l&qa��va����h�u���}�۬�N��g"��dX���N��C�h��	 9G�Ob.�+s���ĩ#؋�X-��k��D��I�㝇_.�
��aϝ�gl6�|V R�������Ԕ ��B��m_?�L��۞k�\ r�C�(؋ClUʘ�迬�;v�w��b`�����C[΋ �+� IhM�@k�����p
W0��_C��bm��<���##´��Yˁ��" �+�̐�@��E���&��/
\B<2�·)�j�|�±�[`�v��J�����2;;��W�-�׋ &�1#s�[Qc�H �S���q:ڟ�74U����oW� �@��g��+a.l�U!��\8�Ï�̔3gP80�[�:1q~�t�H�o��p��q݆�5Cu�O�8ͯ���Żu��gz�"
׼��f<a	�����ƽ¨���.�Q��	W�4'o�K(�j���������(��cm$��MѶz�Dʝ� �>�ѿ	�tVP�����-S ����^6(�Ij˴��VQZ	D�I;EI��P�~���j]�\_*�F,��Ť6�/͜�IPq�	�	�$@�c{RR�2[(@Y �ߙ`��J�"p)�4��i�	*���]>@��A�Tz�*�Y���TL:� ���|O/��O�&�l�;߯Cz���M)����R���� @n}�(�������B��G�q��i[Z�{Y�9���e	�����    IEND�B`� 
BackgroundclWindowNameOpen Workspace (reduced alpha)PngImage.Data
�	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:39+01:00" xmp:ModifyDate="2022-09-01T11:06:02+01:00" xmp:MetadataDate="2022-09-01T11:06:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c87184bb-72dd-4a4b-8017-bd47f89d80f3" xmpMM:DocumentID="adobe:docid:photoshop:eb73ca61-876e-2b4f-a9d1-8143c66bc758" xmpMM:OriginalDocumentID="xmp.did:88a236ff-d429-1e44-b2ab-c5515970910f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:88a236ff-d429-1e44-b2ab-c5515970910f" stEvt:when="2022-06-27T15:59:39+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c87184bb-72dd-4a4b-8017-bd47f89d80f3" stEvt:when="2022-09-01T11:06:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�;�*  �IDATx�Ֆ]L�P�Oal|���h� d%F�1�ɢA��o��|Rj@�AL4Q� EyPc�h0��(N���`p�lk�c�n]��P`=I���m���s�=��@(�̧���A֫O%X�H���o ��7,��R��������BvV��Y9�i��p�h�
p�����p��� ��T�}�3�? dW�9��6@��7�p��k�i) 炾掔�SP]�9�Bk�����K��x��.D���'���%�`. �05�wS t�>�O� �|��}1l���+gR���`_��sf4o���f� �(��HD���\)@;���:�\&@r��(�B����E��9@�e�ig�Y��N-����0n�B¦��	���w ؙ�� :�H�s���ہ���,��CO
��pH�1@xd� ~7(��9�tRFG�F�&(�I=0��p0��#ռݵ��?ֹ��,"rBS|4x]"%N݁�M�#`�� ���`�� =���ȹ{!RF�@H����GU[^���W;0f	����&i���֫HI�@�UU���L��p`T��!8,R�9�qJP"�:S�j}O����4@��S��D�p��	�FƇ���x���:����� ��{�tRF�'P&�&��/��;.��;:4O�@tR��M�-��Jw��n����/ s�������C����@�2hJZ� �n��E�%G-��u�ڭ�1�e?F� ���K����4W��-P���mC)���}KƮ+���k�V�-����G�D �VcN�X|��H�W�0�4���n�6'bBzDDF��z%mX�Ř���fX]R��tCw� �R��x1ƬM#���?�������  ����d/X�    IEND�B`� 
BackgroundclWindowName"Open saved session (reduced alpha)PngImage.Data
�
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:57:55+01:00" xmp:ModifyDate="2022-09-01T10:52:53+01:00" xmp:MetadataDate="2022-09-01T10:52:53+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5fa9d523-f1d1-194c-9f6d-810f3ee83fbc" xmpMM:DocumentID="adobe:docid:photoshop:7fabcb25-b4e0-8e41-ae2d-7f960e61cc87" xmpMM:OriginalDocumentID="xmp.did:b0908b0a-c216-4344-993a-a9e682b0df4e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:b0908b0a-c216-4344-993a-a9e682b0df4e" stEvt:when="2022-06-27T15:57:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5fa9d523-f1d1-194c-9f6d-810f3ee83fbc" stEvt:when="2022-09-01T10:52:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>-�P  _IDATx�ŗklU�����B�T-�]��"��,AmK�D%�1�b�D�|��Z��`���T�(���e�|0b4&��]Ҕ��j�-���8�c3;3��|�&w��w��w�9sf�!"0������� �R�+�C�����������+f����>}�]�9A������걀�~=���Z�2���Q�w�i��׬�mFcC�u�7w�Kg<OjT��`��5�H�� 5o���Oi]?��l����C�v�z�:*�6w�Φ����8~��������MD���x�	�}No���m��]�Y��<�l����ш�ǚ �\.o&�n�ڍN�P�4���:u�z&I���Z��A�j�8�<J��b��B!�^׺���W�F��[��[� T�׀�?=1=��'��jO%z�+-$�2^��!�>�dj "�p�����ٲ*7�V��uho=�0#���n{צxYM(��A�v[�U80��;��وL��/}�9���[�ҖŘ�u�t"(��+�yW�V��Z��X�WliHw?��  ��$'w��X���c���\t�Y��K�ޓGQ���,���Pp%�����@xL� �W�I��oM[ڳQ��U<�Q�,��5;Gut>v2�Ɗ�5��!�-}��2�d������ �����O��Q�&:��y#f7�d�)<߹�[�0ޥ L�0.܎��W)�0О��!�ە����+.���!��j�02��,�C���)72��&XC;C\�}�����%	���g�V�Ȝ���D@2�F�]L�*G�O�1���$��ҨK�V'1�t��PB�=b�gzzb ��q�dЎPz�Z�>I��&�)���?`/��W�N`�K7�N�Dv�Ø���4yt"F��7=�-��>�`��M�F��>�tǌ2�5�G׳�� ��9=�-��ӹ42�Ē��S��J�Fa����}B�?YHLf���|+YJPp~G�����.�Ks�?���ﰔ�f�@W�!4:<C/� �k�G%e�"�f�^�B��1�H��#�6��M���p���3����a��؂aЏ?�5�t �����[i���V�.��5�Q��n8�����d�V�    IEND�B`�  Left�Top�   
TPopupMenuSitesIncrementalSearchPopupMenuLeftTop5 	TMenuItem
MenuItem36ActionSearchSiteNameStartOnlyAction	RadioItem	  	TMenuItem
MenuItem37ActionSearchSiteNameAction	RadioItem	  	TMenuItem
MenuItem38ActionSearchSiteAction	RadioItem	       TPF0TMessageFormMessageFormLeft�Top� BorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionInformationXClientHeight)ClientWidthFColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChanged
TextHeight     TPF0TNonVisualDataModuleNonVisualDataModuleHeight�Widthp TTBXPopupMenuRemoteFilePopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�TopP TTBXItem	TBXItem23ActionCurrentAddEditLinkContextAction  TTBXItemRemoteOpenMenuItemActionCurrentOpenAction  TTBXSubmenuItemRemoteEditMenuItemActionCurrentEditFocusedActionDropdownCombo	OnPopupFocusedEditMenuItemPopup  TTBXSubmenuItemRemoteCopyMenuItemActionRemoteCopyFocusedActionDropdownCombo	 TTBXItem	TBXItem72ActionRemoteCopyFocusedNonQueueAction  TTBXItem	TBXItem69ActionRemoteCopyFocusedQueueAction  TTBXSeparatorItemTBXSeparatorItem9  TTBXItemMoveto1ActionRemoteMoveFocusedAction   TTBXItem
Duplicate3ActionRemoteCopyToFocusedAction  TTBXItemMoveto6ActionRemoteMoveToFocusedAction  TTBXItemDelete1ActionCurrentDeleteFocusedAction  TTBXItemRename1ActionCurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem82Action$CurrentCopyToClipboardFocusedAction2  TTBXSeparatorItemN45  TTBXSubmenuItem!RemoteFilePopupCustomCommandsMenuActionCustomCommandsFileAction TTBXItem    TTBXSubmenuItem
FileNames3Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItemInserttoCommandLine2ActionFileListToCommandLineAction  TTBXItemCopytoClipboard3ActionFileListToClipboardAction  TTBXItemCopytoClipboardIncludePaths3ActionFullFileListToClipboardAction  TTBXItemCopyURLtoClipboard3ActionFileGenerateUrlAction2   TTBXSeparatorItemN1  TTBXItemProperties1ActionCurrentPropertiesFocusedAction   TActionListExplorerActionsImagesGlyphsModule.ExplorerImages	OnExecuteExplorerActionsExecuteOnUpdateExplorerActionsUpdateLeft�Top TActionAutoSizeRemoteColumnsActionTagCategoryColumnsCaption&Automatisk storlekHelpKeywordui_file_panel#widthHint4   Justera kolumnbredden för att passa deras innehållShortCutk@  TActionRemoteCopyQueueActionTagCategoryRemote Selected OperationCaptionLadda ner i &bakgrunden...HelpKeywordtask_downloadHintB   Ladda ner valda fjärrfiler till den lokala katalogen i bakgrunden
ImageIndexk  TActionRemoteCopyFocusedQueueActionTagCategoryRemote Focused OperationCaptionLadda ner i &bakgrunden...HelpKeywordtask_downloadHintB   Ladda ner valda fjärrfiler till den lokala katalogen i bakgrunden
ImageIndexk  TActionLocalCopyQueueActionTag	CategoryLocal Selected OperationCaption   Överför i &bakgrunden...HelpKeywordtask_uploadHint>   Överför valda lokala filer till fjärrkatalogen i bakgrunden
ImageIndexl  TActionLocalCopyFocusedQueueActionTagCategoryLocal Focused OperationCaption   Överför i &bakgrunden...HelpKeywordtask_uploadHint>   Överför valda lokala filer till fjärrkatalogen i bakgrunden
ImageIndexl  TActionRemoteCopyNonQueueActionTagCategoryRemote Selected OperationCaptionLadda &ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionRemoteCopyFocusedNonQueueActionTagCategoryRemote Focused OperationCaptionLadda &ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionLocalCopyNonQueueActionTag	CategoryLocal Selected OperationCaption   &Överför...HelpKeywordtask_uploadHint   Överför|Överför valda filer
ImageIndexX  TActionLocalCopyFocusedNonQueueActionTagCategoryLocal Focused OperationCaption   &Överför...HelpKeywordtask_uploadHint   Överför|Överför valda filer
ImageIndexX  TActionLocalCopyFocusedActionTagCategoryLocal Focused OperationCaption   &Överför...HelpKeywordtask_uploadHint3   Överför|Överför lokala filer till fjärrkatalog
ImageIndexX  TActionRemoteCopyFocusedActionTagCategoryRemote Focused OperationCaption&Ladda ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionRemoteMoveFocusedActionTagCategoryRemote Focused OperationCaptionLadda ner och &ta bort...HelpKeywordtask_downloadHint\   Ladda ner och ta bort|Ladda ner fjärrfiler till den lokala katalogen och ta bort originalet
ImageIndexa  TActionRemoteCopyActionTagCategoryRemote Selected OperationCaptionLadda &ner...HelpKeywordtask_downloadHint9   Ladda ner|Ladda ner fjärrfiler till den lokala katalogen
ImageIndexY  TActionAutoSizeLocalColumnsActionTagCategoryColumnsCaption&Automatisk storlekHelpKeywordui_file_panel#widthHint4   Justera kolumnbredden för att passa deras innehållShortCutk@  TActionResetLayoutRemoteColumnsActionTagCategoryColumnsCaption   Å&terställ layoutHelpKeywordui_file_panel#widthHint;   Återställ till standardlayouten för filpanelens kolumner  TActionGoToTreeActionTagCategoryViewCaption   Gå till trädHelpKeywordui_file_panel#directory_treeHint   Gå till träd
ImageIndexLShortCutT�    TActionLocalTreeActionTagCategoryViewCaption   &TrädHelpKeywordui_file_panel#directory_treeHint   Dölj/visa katalogträd
ImageIndexLShortCutT�    TActionRemoteTreeActionTagCategoryViewCaption   &TrädHelpKeywordui_file_panel#directory_treeHint   Dölj/visa katalogträd
ImageIndexLShortCutT�    TActionQueueItemQueryActionTagCategoryQueueCaption   Vi&sa frågaHelpKeywordui_queue#manageHint'   Visa avvaktande fråga på vald köpost
ImageIndexC  TActionResetLayoutLocalColumnsActionTagCategoryColumnsCaption   Å&terställ layoutHelpKeywordui_file_panel#widthHint;   Återställ till standardlayouten för filpanelens kolumner  TActionQueueItemErrorActionTagCategoryQueueCaption	Vi&sa felHelpKeywordui_queue#manageHint.   Visa avvaktande felmeddelande på vald köpost
ImageIndexD  TActionQueueItemPromptActionTagCategoryQueueCaptionVi&sa promptHelpKeywordui_queue#manageHint'   Visa avvaktande prompt på vald köpost
ImageIndexE  TActionGoToCommandLineActionTagCategoryViewCaption   Gå till komma&ndoradHelpKeywordui_commander#command_lineHint   Gå till kommandoradShortCutM`  TActionQueueItemDeleteActionTagCategoryQueueCaption&AvbrytHelpKeywordui_queue#manageHint   Ta bort vald köpost
ImageIndexG  TActionQueueItemExecuteActionTagCategoryQueueCaption
   &Utför nuHelpKeywordui_queue#manageHintC   Utför vald köpost omedelbart genom att ge den en extra anslutning
ImageIndexF  TActionSelectOneActionTagCategory	SelectionCaption&Markera/avmarkeraHelpKeywordui_file_panel#selecting_filesHint"Markera|Markera/avmarkera vald fil  TActionCurrentRenameActionTagCategorySelected OperationCaption	&Byt namnHelpKeywordtask_renameHint   Byt namn|Byt namn på vald fil
ImageIndex  TActionLocalSortAscendingAction2Tag	CategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintG   Stigande/fallande|Växla stigande/fallande sortering av filer i panelen
ImageIndex%  TActionCurrentEditActionTagCategorySelected OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera markerad fil
ImageIndex9  TActionHideColumnActionTagCategoryColumnsCaption   &Dölj kolumnHelpKeywordui_file_panel#selecting_columnsHint   Dölj kolumn|Dölj vald kolumn  TActionLocalBackActionTag	CategoryLocal DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionRemoteCycleStyleActionTagCategoryStyleCaptionVisaHelpKeywordui_file_panel#view_styleHint9   Visa|Växla mellan att visa olika stilar för katalogvyer
ImageIndex  TActionRemoteIconActionTagCategoryStyleCaptionSt&ora ikonerHelpKeywordui_file_panel#view_styleHintStora ikoner|Visa stora ikoner
ImageIndex  TActionRemoteSmallIconActionTagCategoryStyleCaption   &Små ikonerHelpKeywordui_file_panel#view_styleHint   Små ikoner|Visa små ikoner
ImageIndex	  TActionRemoteListActionTagCategoryStyleCaptionLis&taHelpKeywordui_file_panel#view_styleHintLista|Visa lista
ImageIndex
  TActionRemoteReportActionTagCategoryStyleCaption&Detaljerad listaHelpKeywordui_file_panel#view_styleHint&Detaljerad lista|Visa detaljerad lista
ImageIndex  TActionRemoteMoveToActionTagCategoryRemote Selected OperationCaption&Flytta till...HelpKeywordtask_move_duplicate#moveHint0   Flytta|Flytta markerade filer till fjärrkatalog
ImageIndexd  TActionCurrentDeleteFocusedActionTagCategoryFocused OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesFocusedActionTagCategoryFocused OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionCurrentCreateDirActionTagCategorySelected OperationCaptionS&kapa katalog...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionCurrentDeleteActionTagCategorySelected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionCurrentPropertiesActionTagCategorySelected OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionRemoteBackActionTagCategoryRemote DirectoryCaption	Till&bakaHelpKeywordtask_navigate#special_commands
ImageIndexShortCut%�    TActionRemoteForwardActionTagCategoryRemote DirectoryCaption   &FramåtHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionCommandLinePanelActionTagCategoryViewCaptionKomma&ndoradHelpKeywordui_commander#command_lineHint   Dölj/visa kommandoradShortCutM`  TActionRemoteParentDirActionTagCategoryRemote DirectoryCaption   &Överliggande katalogHelpKeywordtask_navigate#special_commandsHint"   Huvudkatalog|Gå till huvudkatalog
ImageIndexShortCut  TActionRemoteRootDirActionTagCategoryRemote DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHint   Rotkatalog|Gå till rotkatalog
ImageIndexShortCut�@  TActionRemoteHomeDirActionTagCategoryRemote DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHint   Hemkatalog|Gå till hemkatalog
ImageIndex  TActionRemoteRefreshActionTagCategoryRemote DirectoryCaption
&UppdateraHint$   Uppdatera|Uppdatera kataloginnehåll
ImageIndex  TActionAboutActionTagCategoryHelpCaption&Om...HelpKeywordui_aboutHintOm|Visa programinformation
ImageIndexA  TActionStatusBarActionTagCategoryViewCaption   &StatusfältHint   Visa/dölj statusfältet  TActionSessionsTabsAction2TagCategoryViewCaptionFlik&arHint   Visa/dölj flikar  TActionExplorerAddressBandActionTagCategoryViewCaption&AdressHelpKeywordui_toolbarsHint   Visa/dölj adressfältet  TActionExplorerMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHint   Visa/dölj meny  TActionExplorerToolbarBandActionTagCategoryViewCaption&StandardknapparHelpKeywordui_toolbarsHint"   Visa/dölj standardverktygsfältet  TActionRemoteOpenDirActionTagCategoryRemote DirectoryCaption   &Öppna katalog/bokmärkeHelpKeywordtask_navigate#manualHintC   Öppna katalog/bokmärke|Öppna vald katalog eller sparat bokmärke
ImageIndex  TActionSelectActionTagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint Markera|Markera filer efter mask
ImageIndexShortCutk  TActionUnselectActionTagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint$Avmarkera|Avmarkera filer efter mask
ImageIndexShortCutm  TActionSelectAllActionTagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla
ImageIndexShortCutA@  TActionInvertSelectionActionTagCategory	SelectionCaption&Invertera markeringHelpKeywordui_file_panel#selecting_filesHintInvertera markering
ImageIndexShortCutj  TActionExplorerSelectionBandActionTagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för markering  TActionClearSelectionActionTagCategory	SelectionCaption&Rensa markeringHelpKeywordui_file_panel#selecting_filesHintRensa markering
ImageIndexShortCutL`  TActionExplorerSessionBandAction2TagCategoryViewCaptionSessio&ner och flikknapparHelpKeywordui_toolbarsHint4   Dölj/visa verktygsfältet för sessioner och flikar  TActionExplorerPreferencesBandActionTagCategoryViewCaption   InställningsknapparHelpKeywordui_toolbarsHint.   Visa/dölj verktygsfältet för inställningar  TActionExplorerSortBandActionTagCategoryViewCaptionSo&rteringsknapparHelpKeywordui_toolbarsHint)   Visa/dölj verktygsfältet för sortering  TActionExplorerUpdatesBandActionTagCategoryViewCaption&UppdateringsknappHelpKeywordui_toolbarsHint+   Dölj/visa verktygsfält för uppdateringar  TActionExplorerTransferBandActionTagCategoryViewCaption   &Överför inställningarHelpKeywordui_toolbarsHint9   Dölj/visa verktygsfält för överföringsinställningar  TAction ExplorerCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionSiteManagerActionTagCategorySessionCaption&Hantera webbplats...HelpKeywordui_loginHints   Hantera webbplats|Öppnar hantera webbplats (håll ner Shift för att öppna hantera webbplats i ett nytt fönster)  TActionCloseTabActionTagCategoryTabCaption   &Stäng flikHelpKeywordui_tabs#workingHint   Stäng den aktuella fliken
ImageIndexSecondaryShortCuts.StringsCtrl+W ShortCutD`  TActionDisconnectSessionActionTagCategorySessionCaption   &Koppla ifrån sessionHelpKeywordtask_connections#closingHint=   Koppla ifrån den aktuella sessionen, men håll fliken öppen
ImageIndext  TActionReconnectSessionActionTagCategorySessionCaption   Å&teranslut sessionHelpKeywordtask_connectionsHint0   Återanslut den aktuella frånkopplade sessionenShortCutR`  TActionSavedSessionsAction2TagCategorySessionCaptionWebb&platserHelpKeyword.task_connections#opening_additional_connectionHint   Öppna webbplats
ImageIndex  TActionWorkspacesActionTagCategoryTabCaption&ArbetsytorHelpKeyword	workspaceHint   Öppna arbetsyta
ImageIndexe  TActionPreferencesActionTagCategoryViewCaption   &Inställningar...HelpKeywordui_preferencesHint2   Inställningar|Visa/ändra användarinställningar
ImageIndexShortCutP�    TActionRemoteChangePathAction2TagCategoryRemote DirectoryCaption&Byt katalogHelpKeywordtask_navigateHint-   Tillåter val av olika kataloger för panelen
ImageIndexShortCutq�    TActionLocalForwardActionTag	CategoryLocal DirectoryCaption   &FramåtHelpKeywordtask_navigate#special_commands
ImageIndexShortCut'�    TActionLocalParentDirActionTagCategoryLocal DirectoryCaption&HuvudkatalogHelpKeywordtask_navigate#special_commandsHint"   Huvudkatalog|Gå till huvudkatalog
ImageIndexShortCut  TActionLocalRootDirActionTagCategoryLocal DirectoryCaption&RotkatalogHelpKeywordtask_navigate#special_commandsHint    Rotkatalog|Gå till rotkatalogen
ImageIndexShortCut�@  TActionLocalHomeDirActionTag	CategoryLocal DirectoryCaption&HemkatalogHelpKeywordtask_navigate#special_commandsHint    Hemkatalog|Gå till hemkatalogen
ImageIndex  TActionLocalRefreshActionTag	CategoryLocal DirectoryCaption
&UppdateraHint$   Uppdatera|Uppdatera kataloginnehåll
ImageIndex  TActionLocalOpenDirActionTag	CategoryLocal DirectoryCaption   &Öppna katalog/bokmärke...HelpKeywordtask_navigate#manualHintC   Öppna katalog/bokmärke|Öppna vald katalog eller sparat bokmärke
ImageIndex  TActionLocalChangePathAction2TagCategoryLocal DirectoryCaption
&Byt enhetHelpKeywordtask_navigateHint)   Tillåter val av olika enheter för panel
ImageIndexShortCutp�    TActionToolBar2ActionTagCategoryViewCaption   Verktygsfält snabb&tangenterHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för snabbtangenter  TActionCommanderMenuBandActionTagCategoryViewCaption&MenyHelpKeywordui_toolbarsHint   Dölj/visa meny  TActionCommanderSessionBandAction2TagCategoryViewCaptionSessio&ner och flikknapparHelpKeywordui_toolbarsHint4   Dölj/visa verktygsfältet för sessioner och flikar  TActionCommanderPreferencesBandActionTagCategoryViewCaption   InställningsknapparHelpKeywordui_toolbarsHint.   Dölj/visa verktygsfältet för inställningar  TActionCommanderSortBandActionTagCategoryViewCaptionS&orteringsknapparHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfältet för sortering  TActionCommanderUpdatesBandActionTagCategoryViewCaption&UppdateringsknappHelpKeywordui_toolbarsHint)   Dölj/visa verktygsfält för uppdatering  TActionCommanderTransferBandActionTagCategoryViewCaption   ÖverföringsinställningarHelpKeywordui_toolbarsHint9   Dölj/visa verktygsfält för överföringsinställningar  TActionCommanderCommandsBandActionTagCategoryViewCaption&KommandoknapparHelpKeywordui_toolbarsHint)   Visa/dölj verktygsfältet för kommandon  TAction!CommanderCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TAction CommanderLocalHistoryBandAction2TagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint#   Dölj/visa verktygsfältet historik  TAction#CommanderLocalNavigationBandAction2TagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint%   Dölj/visa verktygsfältet navigering  TActionCommanderLocalFileBandAction2TagCategoryViewCaption&FilknapparHelpKeywordui_toolbarsHint   Dölj/visa verktygsfältet fil  TAction"CommanderLocalSelectionBandAction2TagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint$   Dölj/visa verktygsfältet markering  TAction!CommanderRemoteHistoryBandAction2TagCategoryViewCaption&HistorikknapparHelpKeywordui_toolbarsHint#   Dölj/visa verktygsfältet historik  TAction$CommanderRemoteNavigationBandAction2TagCategoryViewCaption&NavigeringsknapparHelpKeywordui_toolbarsHint%   Dölj/visa verktygsfältet navigering  TActionCommanderRemoteFileBandAction2TagCategoryViewCaption&FilknapparHelpKeywordui_toolbarsHint   Dölj/visa verktygsfältet fil  TAction#CommanderRemoteSelectionBandAction2TagCategoryViewCaption&MarkeringsknapparHelpKeywordui_toolbarsHint$   Dölj/visa verktygsfältet markering  TActionLocalStatusBarAction2TagCategoryViewCaption   Statusf&ältHint   Dölj/visa panelens statusfält  TActionRemoteStatusBarAction2TagCategoryViewCaption   Statusf&ältHint   Dölj/visa panelens statusfält  TActionLocalSortByNameAction2Tag	CategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint+Sortera efter namn|Sortera panel efter namn
ImageIndexShortCutr@  TActionLocalSortByExtAction2Tag	CategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHint9   Sortera efter filändelse|Sortera panel efter filändelse
ImageIndex ShortCuts@  TActionLocalSortBySizeAction2Tag	CategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint4Sortera efter storlek|Sortera panel efter filstorlek
ImageIndex#ShortCutu@  TActionLocalSortByAttrAction2Tag	CategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHint3Sortera efter attribut|Sortera panel efter attribut
ImageIndex$ShortCutv@  TActionLocalSortByTypeAction2Tag	CategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint,Sortera efter typ|Sortera panel efter filtyp
ImageIndex"  TActionLocalSortByChangedAction2Tag	CategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHint:   Sortera efter tid|Sortera panel efter senaste ändringstid
ImageIndex!ShortCutt@  TActionRemoteSortAscendingAction2TagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintG   Stigande/fallande|Växla stigande/fallande sortering av filer i panelen
ImageIndex%  TActionRemoteSortByNameAction2TagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint+Sortera efter namn|Sortera panel efter namn
ImageIndexShortCutr@  TActionRemoteSortByExtAction2TagCategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHint9   Sortera efter filändelse|Sortera panel efter filändelse
ImageIndex ShortCuts@  TActionRemoteSortBySizeAction2TagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint4Sortera efter storlek|Sortera panel efter filstorlek
ImageIndex#ShortCutu@  TActionRemoteSortByRightsAction2TagCategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHint3Sortera efter attribut|Sortera panel efter attribut
ImageIndex$ShortCutv@  TActionRemoteSortByChangedAction2TagCategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHint:   Sortera efter tid|Sortera panel efter senaste ändringstid
ImageIndex!ShortCutt@  TActionRemoteSortByOwnerAction2TagCategorySortCaption   Efter ä&gareHelpKeywordui_file_panel#sorting_filesHint2   Sortera efter ägare|Sortera panel efter filägare
ImageIndex&ShortCutw@  TActionRemoteSortByGroupAction2TagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHint0Sortera efter grupp|Sortera panel efter filgrupp
ImageIndex'ShortCutx@  TActionRemoteSortByTypeAction2TagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint,Sortera efter typ|Sortera panel efter filtyp
ImageIndex"  TActionCurrentSortAscendingActionTagCategorySortCaption	Stig&andeHelpKeywordui_file_panel#sorting_filesHintW   Stigande/fallande|Växla sortering mellan stigande och fallande ordning i aktuell panel
ImageIndex%  TActionCurrentSortByNameActionTagCategorySortCaptionEfter &namnHelpKeywordui_file_panel#sorting_filesHint3Sortera efter namn|Sortera aktuell panel efter namn
ImageIndexShortCutr@  TActionCurrentSortByExtActionTagCategorySortCaption   Efter &filändelseHelpKeywordui_file_panel#sorting_filesHintA   Sortera efter filändelse|Sortera aktuell panel efter filändelse
ImageIndex ShortCuts@  TActionCurrentSortBySizeActionTagCategorySortCaptionEfter &storlekHelpKeywordui_file_panel#sorting_filesHint<Sortera efter storlek|Sortera aktuell panel efter filstorlek
ImageIndex#ShortCutu@  TActionCurrentSortByTypeAction2TagCategorySortCaptionEfter fil&typHelpKeywordui_file_panel#sorting_filesHint4Sortera efter typ|Sortera aktuell panel efter filtyp
ImageIndex"  TActionCurrentSortByRightsActionTagCategorySortCaptionEfter &attributHelpKeywordui_file_panel#sorting_filesHintK   Sortera efter attribut|Sortera aktuell panel efter attribut/filrättigheter
ImageIndex$ShortCutv@  TActionCurrentSortByChangedActionTagCategorySortCaption   Efter senast &ändradHelpKeywordui_file_panel#sorting_filesHintH   Sortera efter senast &ändrad|Sortera aktuell panel efter senast ändrad
ImageIndex!ShortCutt@  TActionCurrentSortByOwnerActionTagCategorySortCaption   Efter ä&gareHelpKeywordui_file_panel#sorting_filesHintO   Sortera efter ägare|Sortera aktuell panel efter filägare (endast fjärrpanel)
ImageIndex&ShortCutw@  TActionCurrentSortByGroupActionTagCategorySortCaptionEfter &gruppHelpKeywordui_file_panel#sorting_filesHintM   Sortera efter grupp|Sortera fjärrpanelen efter filgrupp (endast fjärrpanel)
ImageIndex'ShortCutx@  TActionSortColumnAscendingActionTagCategorySortCaptionSortera stig&andeHelpKeywordui_file_panel#sorting_filesHint(Sortera filer stigande efter vald kolumn
ImageIndex)  TActionSortColumnDescendingActionTagCategorySortCaptionSortera fallan&deHelpKeywordui_file_panel#sorting_filesHint(Sortera filer fallande efter vald kolumn
ImageIndex(  TActionHomepageActionTagCategoryHelpCaptionProdukt&hemsidaHint9   Öppnar webbläsaren och går till applikationens hemsida
ImageIndex*  TActionHistoryPageActionTagCategoryHelpCaption&VersionshistorikHintO   Öppnar webbläsaren och går till webbsida med applikationens versionshistorik  TActionSaveCurrentSessionAction2TagCategorySessionCaption&Spara session som webbplats...HelpKeywordtask_connections#savingHint?Spara session som webbplats|Spara aktuell session som webbplats
ImageIndex+  TActionShowHideRemoteNameColumnAction2TagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen namn
ImageIndex,  TActionShowHideRemoteExtColumnAction2TagCategoryColumnsCaption   &FiländelseHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen filändelse
ImageIndex-  TActionShowHideRemoteSizeColumnAction2TagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen storlek
ImageIndex/  TAction"ShowHideRemoteChangedColumnAction2TagCategoryColumnsCaption   Se&nast ändradHelpKeywordui_file_panel#selecting_columnsHint"   Visa/dölj kolumnen senast ändrad
ImageIndex0  TAction!ShowHideRemoteRightsColumnAction2TagCategoryColumnsCaption   Fil&rättigheterHelpKeywordui_file_panel#selecting_columnsHint#   Visa/dölj kolumnen filrättigheter
ImageIndex1  TAction ShowHideRemoteOwnerColumnAction2TagCategoryColumnsCaption   &ÄgareHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen ägare
ImageIndex2  TAction ShowHideRemoteGroupColumnAction2TagCategoryColumnsCaption&GruppHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen grupp
ImageIndex3  TAction%ShowHideRemoteLinkTargetColumnAction2TagCategoryColumnsCaption
   &LänkmålHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen länkmål
ImageIndexR  TActionShowHideRemoteTypeColumnAction2TagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen filtyp
ImageIndex.  TActionShowHideLocalNameColumnAction2TagCategoryColumnsCaption&NamnHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen namn
ImageIndex,  TActionShowHideLocalExtColumnAction2TagCategoryColumnsCaption   &FiländelseHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen filändelse
ImageIndex-  TActionShowHideLocalTypeColumnAction2TagCategoryColumnsCaptionFil&typHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen filtyp
ImageIndex.  TActionShowHideLocalSizeColumnAction2TagCategoryColumnsCaption&StorlekHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen storlek
ImageIndex/  TAction!ShowHideLocalChangedColumnAction2TagCategoryColumnsCaption   Senast &ändradHelpKeywordui_file_panel#selecting_columnsHint"   Visa/dölj kolumnen senast ändrad
ImageIndex0  TActionShowHideLocalAttrColumnAction2TagCategoryColumnsCaption	&AttributHelpKeywordui_file_panel#selecting_columnsHint   Visa/dölj kolumnen attribut
ImageIndex1  TActionCompareDirectoriesAction2TagCategoryCommandCaption   &Jämför katalogerHelpKeywordtask_compare_directoriesHint8   Jämför kataloger|Markera olika filer mellan filpaneler
ImageIndex4ShortCutq   TActionSynchronizeActionTagCategoryCommandCaption!   &Håll fjärrkatalogen uppdateradHelpKeywordtask_keep_up_to_dateHintA   Håll fjärrkatalogen uppdaterad|Håll fjärrkatalogen uppdaterad
ImageIndex5ShortCutU@  TActionForumPageActionTagCategoryHelpCaption&SupportforumHint=   Öppnar webbläsaren och gå till webbsida med supportforumet  TActionLocalAddBookmarkAction2Tag	CategoryLocal DirectoryCaption   &Lägg till bokmärkenHelpKeywordtask_navigate#bookmarksHintL   Lägg till i bokmärken|Lägg till den aktuella katalogen i bokmärkeslistan
ImageIndex6ShortCutB@  TActionRemoteAddBookmarkAction2TagCategoryRemote DirectoryCaption   &Lägg till bokmärkenHelpKeywordtask_navigate#bookmarksHintL   Lägg till i bokmärken|Lägg till den aktuella katalogen i bokmärkeslistan
ImageIndex6ShortCutB@  TActionConsoleActionTagCategoryCommandCaption   Öppna &terminalfönsterHelpKeyword
ui_consoleHint�   Öppna terminalfönster|Öppnar terminalfönster som tillåter körande av godtyckligt extrakommando (med undantag av de som kräver användarinput)
ImageIndex7ShortCutT`  TActionPuttyActionTagCategoryCommandCaption   Öppna session i &PuTTYHelpKeywordintegration_putty#open_puttyHintZ   Öppna session i PuTTY|Starta PuTTY SSH-terminalprogram och öppna aktuell session med den
ImageIndex@ShortCutP@  TActionLocalExploreDirectoryActionTag	CategoryLocal DirectoryCaption&Utforska katalogHint+   Öppnar utforskaren i aktuell lokal katalog
ImageIndex8ShortCutE�    TActionCurrentOpenActionTagCategoryFocused OperationCaption   &ÖppnaHelpKeyword	task_editHintQ   Öppna dokument|Öppnar valt dokument med program som filtypen är associerad med
ImageIndex:  TActionSynchronizeBrowsingAction2TagCategoryCommand	AutoCheck	Caption   Synkronisera &bläddringHelpKeyword"task_navigate#synchronize_browsingHintF   Synkronisera bläddring|Synkronisera bläddring mellan båda panelerna
ImageIndex;ShortCutB�    TActionCurrentAddEditLinkActionTagCategorySelected OperationCaption   Lägg till/redigera &länk...HelpKeyword	task_linkHintZ   Lägg till/redigera länk|Lägger till ny länk/genväg eller redigerar vald länk/genväg
ImageIndex<  TActionCurrentAddEditLinkContextActionTagCategorySelected OperationCaption   Redigera &länk...HelpKeyword	task_linkHint*   Redigera länk|Redigera vald länk/genväg
ImageIndex<  TActionCloseApplicationAction2TagCategoryCommandCaption&AvslutaHintH   Avsluta applikation|Stäng applikation (alla öppnade sessioner stängs)
ImageIndex=  TActionOpenedTabsActionTagCategoryTabCaption   Ö&ppna flikarHelpKeywordui_tabs#switchHint'   Välj flik|Välj flik för att aktivera
ImageIndex>  TActionDuplicateTabActionTagCategoryTabCaptionDu&plicera flikHelpKeywordui_tabsHinte   Duplicera flik|Öppna ny flik med samma mapp (håll ned Skift för att öppna fliken i nytt fönster)
ImageIndex[  TActionNewLinkActionTagCategoryCommandCaption	   &Länk...HelpKeyword	task_linkHint"   Skapa länk|Skapa ny länk/genväg
ImageIndex<  TActionCustomCommandsFileActionTagCategoryCommandCaptionFiler &anpassade kommandonHelpKeywordcustom_commandHint%   Kör anpassade kommandon på vald fil  TActionCustomCommandsNonFileActionTagCategoryCommandCaptionStatiska &anpassade kommandonHelpKeywordcustom_commandHint4   Kör anpassade kommandon som inte fungerar på filer  TActionCustomCommandsCustomizeActionTagCategoryCommandCaption&Anpassa...HelpKeywordui_pref_commandsHintAnpassa egna kommandon
ImageIndex  TActionCustomCommandsEnterActionTagCategoryCommandCaption   Lä&gg in...HelpKeyword(custom_command#executing_and_configuringHint#   Lägg in egna kommandon för ad hoc
ImageIndexZ  TAction CustomCommandsEnterFocusedActionTagCategoryCommandCaption   Lä&gg in...HelpKeyword(custom_command#executing_and_configuringHint#   Lägg in egna kommandon för ad hoc
ImageIndexZ  TActionCheckForUpdatesActionTagCategoryHelpCaption   Sök efter &uppdateringarHelpKeywordupdatesHint0   Frågar applikationens webbsida om uppdateringar
ImageIndex?  TActionDonatePageActionTagCategoryHelpCaption&DoneraHintG   Öppnar webbläsaren och går till programmets webbsida för donationer  TActionCustomCommandsLastActionTagCategoryCommandCaptionCustomCommandsLastActionHelpKeyword(custom_command#executing_and_configuring  TActionCustomCommandsLastFocusedActionTagCategoryCommandCaptionCustomCommandsLastFocusedActionHelpKeyword(custom_command#executing_and_configuring  TActionFileSystemInfoActionTagCategoryCommandCaption&Server/protokollinformationHelpKeyword	ui_fsinfoHint Visa server/protokollinformation
ImageIndex  TActionClearCachesActionTagCategoryCommandCaption&Rensa cacheHelpKeyworddirectory_cacheHint1   Rensa cache för kataloglistning och katalogbyten  TActionFullSynchronizeActionTagCategoryCommandCaption&Synkronisera...HelpKeywordtask_synchronize_fullHint,   Synkronisera lokal katalog med fjärrkatalog
ImageIndexBShortCutS@  TActionRemoteMoveToFocusedActionTagCategoryRemote Focused OperationCaption&Flytta till...HelpKeywordtask_move_duplicate#moveHint0   Flytta|Flytta markerade filer till fjärrkatalog
ImageIndexd  TActionShowHiddenFilesActionTagCategoryViewCaption   Visa/dölj &dolda filerHelpKeywordui_file_panel#hidden_filesHint)   Växla visning av dolda filer i panel(er)ShortCutH�    TActionFormatSizeBytesNoneActionTagCategoryViewCaption&ByteHelpKeywordui_pref_panels#commonHintVisa filstorlekar i byte  TActionLocalPathToClipboardAction2TagCategoryLocal DirectoryCaption   Kopiera s&ökväg till urklippHelpKeywordfilenames#cwdHint,   Kopiera den aktuella sökvägen till urklipp  TActionRemotePathToClipboardAction2TagCategoryRemote DirectoryCaption   Kopiera s&ökväg till urklippHelpKeywordfilenames#cwdHint,   Kopiera den aktuella sökvägen till urklipp  TActionFileListToCommandLineActionTagCategorySelected OperationCaptionIn&foga till kommandoradHelpKeywordfilenames#command_lineHint/Infoga markerade filers namn till kommandoradenShortCut@  TActionFileListToClipboardActionTagCategorySelected OperationCaption&Kopiera till urklippHelpKeywordfilenames#file_nameHint*Kopiera markerade filers namn till urklippShortCutC`  TActionFullFileListToClipboardActionTagCategorySelected OperationCaption,   Kopiera till urklipp (inklusive s&ökvägar)HelpKeywordfilenames#file_nameHint=   Kopiera markerade filers namn inklusive sökväg till urklippShortCutC�    TActionQueueGoToActionTagCategoryQueueCaption	   &Gå tillHelpKeywordui_queue#manageHint   Gå till överföringskölistan
ImageIndexJShortCutQ@  TActionQueueItemUpActionTagCategoryQueueCaptionFlytta &uppHelpKeywordui_queue#manageHint2   Flytta upp vald köpost för att utföras tidigare
ImageIndexH  TActionQueueItemDownActionTagCategoryQueueCaptionFlytta &nerHelpKeywordui_queue#manageHint0   Flytta ner vald köpost för att utföras senare
ImageIndexI  TActionQueueToggleShowActionTagCategoryQueueCaption   &KöHint   Visa/dölj kölista
ImageIndexJ  TActionQueueShowActionTagCategoryQueueCaptionVi&saHelpKeywordui_queueHint   Visa kölista  TActionQueueHideWhenEmptyActionTagCategoryQueueCaption   Dölj ifall &tomHelpKeywordui_queueHint    Dölj kölistan när den är tom  TActionQueueHideActionTagCategoryQueueCaption   &DöljHelpKeywordui_queueHint   Dölj kölista  TActionQueueToolbarActionTagCategoryQueueCaption   &VerktygsfältHint@   Dölj/visa verktygsfältet för kölistan (på kölistans panel)  TActionQueueFileListActionTagCategoryQueueCaption	&FillistaHint#   Dölj/visa fullständig köfillista  TActionQueueResetLayoutColumnsActionTagCategoryQueueCaption   Å&terställ kolumnlayoutHint3   Återställ till standardlayouten för listkolumner  TActionQueuePreferencesActionTagCategoryQueueCaptionA&npassa...HelpKeywordui_pref_backgroundHint   Anpassa kölista
ImageIndex  TActionPasteAction3TagCategoryCommandCaption   &Klistra in från urklippHelpKeyword	clipboardHint�   Klistra in filer från urklipp till aktuell katalog i aktiv panel; eller öppnar sökväg från urklipp i aktiv panel; eller öppnar sessions-URL från urklipp
ImageIndexKShortCutV@  TActionNewFileActionTagCategoryCommandCaption&Fil...HelpKeyword	task_editHint1   Skapa fil|Skapar ny fil och öppnas den i editorn
ImageIndexM  TActionEditorListCustomizeActionTagCategoryCommandCaption&Konfigurera...HelpKeywordui_pref_editorHint   Skräddarsy editorer
ImageIndex  TActionRemoteCopyToFocusedActionTagCategoryRemote Focused OperationCaption&Dubblera...HelpKeywordtask_move_duplicate#duplicateHint3   Dubblera|Dubbleras valda filer till fjärrkatalogen
ImageIndexN  TActionRemoteCopyToActionTagCategoryRemote Selected OperationCaption&Dubblera...HelpKeywordtask_move_duplicate#duplicateHint2   Dubblera|Dubblera valda filer till fjärrkatalogen
ImageIndexN  TActionFileGenerateUrlAction2TagCategorySelected OperationCaptionSkapa fil-&URL...HelpKeywordui_generateurlHint   Skapa URL:er för valda filer  TActionTableOfContentsActionTagCategoryHelpCaption
   I&nnehållHintI   Öppnar webbläsare och går till dokumentationens innehållsförteckning
ImageIndexOShortCutp  TActionFileListFromClipboardActionTagCategorySelected OperationCaption&Transfer Files in ClipboardHelpKeyword	clipboardHint+Transfer files whose names are in clipboard  TActionLocalCopyActionTag	CategoryLocal Selected OperationCaption   &Överför...HelpKeywordtask_uploadHint   Överför|Överför valda filer
ImageIndexX  TActionCurrentDeleteAlternativeActionTagCategorySelected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort valda filer
ImageIndex  TActionCurrentEditWithActionTagCategorySelected OperationCaptionRedigera &med...HelpKeyword	task_editHint9Redigera med|Redigera valda filer med editorn som ni valt  TActionDownloadPageActionTagCategoryHelpCaption
Ladda &nerHintA   Öppnar webbläsare och går till applikationens nerladdningssida  TActionUpdatesPreferencesActionTagCategoryHelpCaptionKonfi&gurera...HelpKeywordui_pref_updatesHintC   Konfigurera automatisk kontroll av uppdateringar för applikationen
ImageIndex  TActionFormatSizeBytesKilobytesActionTagCategoryViewCaption	&KilobyteHelpKeywordui_pref_panels#commonHintVisa filstorlekar i kilobyte  TActionFormatSizeBytesShortActionTagCategoryViewCaption&Kort formatHelpKeywordui_pref_panels#commonHintVisa filstorlekar i kort format  TActionPresetsPreferencesActionTagCategoryViewCaption&Konfigurera...HelpKeywordui_pref_transferHint2   Konfigurera förinställningar för överföringar
ImageIndex  TActionLockToolbarsActionTagCategoryViewCaption   &Lås verktygsfältHelpKeywordui_toolbarsHint3   Hindra flyttning och dockning av alla verktygsfält  TActionSelectiveToolbarTextActionTagCategoryViewCaption&Visa valbara textetiketterHelpKeywordui_toolbarsHintD   Visa textetiketter på utvalda viktiga kommandon på verktygsfältet  TActionToolbarIconSizeActionTagCategoryViewCaption!   St&orlek på verktygsfältsikonerHelpKeywordui_toolbarsHint'   Ändra storlek på verktygsfältsikoner  TActionToolbarIconSizeNormalActionTagCategoryViewCaption&NormalHelpKeywordui_toolbarsHint!   Visa normala verktygsfältsikoner  TActionToolbarIconSizeLargeActionTagCategoryViewCaption&StoraHelpKeywordui_toolbarsHint   Visa stora verktygsfältsikoner  TActionToolbarIconSizeVeryLargeActionTagCategoryViewCaption&Mycket storaHelpKeywordui_toolbarsHint&   Visa mycket stora verktygsfältsikoner  TActionCustomCommandsBandActionTagCategoryViewCaptionEgna ko&mmandoknapparHelpKeywordui_toolbarsHint,   Dölj/visa verktygsfält för egna kommandon  TActionColorMenuAction2TagCategoryViewCaption   F&ärgHelpKeywordtask_connections#session_colorHint$   Ändra färg på den aktuella fliken  TActionAutoReadDirectoryAfterOpActionTagCategoryViewCaptionLadda auto&matisk om katalogHint=   Ändra automatisk omladdning av fjärrkatalog efter operationShortCutR�    TActionQueueItemPauseActionTagCategoryQueueCaption&PausaHelpKeywordui_queue#manageHint   Pausa vald köpost
ImageIndexS  TActionQueueItemResumeActionTagCategoryQueueCaption   &ÅterupptaHelpKeywordui_queue#manageHint   Återuppta vald pausad köpost
ImageIndexF  TActionQueuePauseAllActionTagCategoryQueueCaption&Pausa allaHelpKeywordui_queue#manageHint   Pausa alla köposter som körs
ImageIndexT  TActionQueueResumeAllActionTagCategoryQueueCaption   &Återuppta allaHelpKeywordui_queue#manageHint!   Återuppta alla pausade köposter
ImageIndexU  TActionQueueDeleteAllDoneActionTagCategoryQueueCaption   Ta bort alla &slutfördaHelpKeywordui_queue#manageHint!   Ta bort alla slutförda köposter
ImageIndexc  TActionQueueEnableActionTagCategoryQueueCaption   &ProcessköHelpKeywordui_queue#manageHints   Aktivera köbehandling|Aktivera köbehandling (väntande köposter startar inte, när köbehandling är inaktiverad
ImageIndex`ShortCutQ`  TActionQueueDisconnectOnceEmptyAction2TagCategoryQueueCaption   &Koppla ifrån sessionHelpKeywordui_queueHint'   Koppla ifrån session när kön är tom
ImageIndexW  TActionRestoreSelectionActionTagCategory	SelectionCaption   &Återställ markeringHelpKeywordui_file_panel#selecting_filesHint"   Återställ föregående markering
ImageIndexVShortCutS`  TActionLocalSelectAction2TagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint Markera|Markera filer efter mask
ImageIndex  TActionLocalUnselectAction2TagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint$Avmarkera|Avmarkera filer efter mask
ImageIndex  TActionLocalSelectAllAction2TagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla
ImageIndex  TActionCurrentEditFocusedActionTagCategoryFocused OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera valda filer
ImageIndex9  TActionCurrentEditWithFocusedActionTagCategoryFocused OperationCaptionRedigera &med...HelpKeyword	task_editHint9Redigera med|Redigera valda filer med editorn som ni valt  TActionNewDirActionTagCategoryCommandCaptionKatalo&g...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionQueueShutDownOnceEmptyAction2TagCategoryQueueCaption   Stäng av datornHelpKeywordui_queueHint"   Stäng av datorn när kön är tom
ImageIndex]  TActionQueueSuspendOnceEmptyAction2TagCategoryQueueCaption   Försätt datorn i vilolägeHelpKeywordui_queueHint.   Försätt datorn i viloläge när kön är tom
ImageIndexi  TActionQueueIdleOnceEmptyActionTagCategoryQueueCaption   &Förbli inaktivChecked	HelpKeywordui_queueHint!   Förbli inaktiv när kön är tom
ImageIndex^  TActionQueueCycleOnceEmptyActionTagCategoryQueueCaption   &Tom köHelpKeywordui_queueHint1   Ändra åtgärd som ska utföras då kön är tom
ImageIndex^  TTBEditActionQueueItemSpeedActionTagCategoryQueueHelpKeywordui_queue#manageHint)   Ändra hastighetsgräns för vald köpost
ImageIndexmEditCaption
&Hastighet  TActionQueueDeleteAllActionTagCategoryQueueCaption&Avbryt allaHelpKeywordui_queue#manageHint   Ta bort alla köposter
ImageIndexj  TActionLocalFilterActionTag	CategoryLocal DirectoryCaption&Filtrera...HelpKeywordui_file_panel#filteringHintFiltrera|Filtrera visade filer
ImageIndex\ShortCutF�    TActionRemoteFilterActionTagCategoryRemote DirectoryCaption
&Filter...HelpKeywordui_file_panel#filteringHintFilter|Filtrera visade filer
ImageIndex\ShortCutF�    TActionRemoteFindFilesAction2TagCategoryRemote DirectoryCaption   Sö&k filer..HelpKeyword	task_findHint%Hitta filer|Hitta filer och kataloger
ImageIndex_  TActionCurrentEditInternalActionTagCategorySelected OperationCaption&Intern editorHelpKeyword	task_editHint8Redigera (intern)|Redigera valda filer med intern editor  TActionSaveWorkspaceActionTagCategoryTabCaptionSpara arbets&yta...HelpKeyword	workspaceHintSpara arbetsyta|Spara arbetsyta
ImageIndexf  TActionLocalRenameAction2TagCategoryLocal Selected OperationCaption	&Byt namnHelpKeywordtask_renameHint   Byt namn|Byt namn på vald fil
ImageIndex  TActionLocalEditAction2TagCategoryLocal Selected OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera markerad fil
ImageIndex9  TActionLocalMoveActionTag	CategoryLocal Selected OperationCaption   Överför och ta &bort...HelpKeywordtask_uploadHint]   Överför och ta bort|Överför valda lokala filer till fjärrkatalogen och tar bort original
ImageIndexb  TActionLocalCreateDirAction3TagCategoryLocal Selected OperationCaptionKatalo&g...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionLocalDeleteAction2TagCategoryLocal Selected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionLocalPropertiesAction2TagCategoryLocal Selected OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionLocalAddEditLinkAction3TagCategoryLocal Selected OperationCaption   &Genväg...HelpKeyword	task_linkHintZ   Lägg till/redigera länk|Lägger till ny länk/genväg eller redigerar vald länk/genväg
ImageIndex<  TActionRemoteRenameAction2TagCategoryRemote Selected OperationCaption	&Byt namnHelpKeywordtask_renameHint   Byt namn|Byt namn på vald fil
ImageIndex  TActionRemoteEditAction2TagCategoryRemote Selected OperationCaption	&RedigeraHelpKeyword	task_editHintRedigera|Redigera markerad fil
ImageIndex9  TActionRemoteMoveActionTagCategoryRemote Selected OperationCaptionLadda ner och &ta bortHelpKeywordtask_downloadHintY   Ladda ner och ta bort|Ladda ner valda fjärrfiler till lokal katalog och ta bort original
ImageIndexa  TActionRemoteCreateDirAction3TagCategoryRemote Selected OperationCaptionKatalo&g...HelpKeywordtask_create_directoryHintSkapa katalog|Skapa ny katalog
ImageIndex  TActionRemoteDeleteAction2TagCategoryRemote Selected OperationCaption&Ta bortHelpKeywordtask_deleteHintTa bort|Ta bort markerade filer
ImageIndex  TActionRemotePropertiesAction2TagCategoryRemote Selected OperationCaption&EgenskaperHelpKeywordtask_propertiesHint6   Egenskaper|Visa/ändra egenskaper för markerade filer
ImageIndex  TActionRemoteAddEditLinkAction3TagCategoryRemote Selected OperationCaption	   &Länk...HelpKeyword	task_linkHintZ   Lägg till/redigera länk|Lägger till ny länk/genväg eller redigerar vald länk/genväg
ImageIndex<  TActionRemoteSelectAction2TagCategory	SelectionCaption&Markera filerHelpKeyword	ui_selectHint Markera|Markera filer efter mask
ImageIndex  TActionRemoteUnselectAction2TagCategory	SelectionCaptionA&vmarkera filerHelpKeyword	ui_selectHint$Avmarkera|Avmarkera filer efter mask
ImageIndex  TActionRemoteSelectAllAction2TagCategory	SelectionCaptionM&arkera allaHelpKeywordui_file_panel#selecting_filesHintMarkera alla
ImageIndex  TActionLocalMoveFocusedActionTagCategoryLocal Focused OperationCaption   Överför och &ta bort...HelpKeywordtask_uploadHintZ   Överför och ta bort|Överför valda lokala filer till fjärrkatalog och ta bort original
ImageIndexb  TAction CurrentEditInternalFocusedActionTagCategoryFocused OperationCaption&Intern editorHelpKeyword	task_editHint8Redigera (intern)|Redigera valda filer med intern editor  TActionCurrentSystemMenuFocusedActionTagCategoryFocused OperationCaption&SystemmenyHintn   Visa filsystemets snabbmeny (i egenskaper kan du välja att visa den som standard istället för inbyggd meny)  TActionSessionGenerateUrlAction2TagCategorySessionCaptionSkapa sessions-&URL/kod...HelpKeywordui_generateurlHint/   Skapa URL eller kod för den aktuella sessionen  TActionSelectSameExtActionTagCategory	SelectionCaption$   &Markera filer med samma filtilläggHint:   Markera alla filer med samma filtillägg som fokuserad filShortCutk�    TActionUnselectSameExtActionTagCategory	SelectionCaption&   &Avmarkera filer med samma filtilläggHint<   Avmarkera alla filer med samma filtillägg som fokuserad filShortCutm�    TActionGoToAddressActionTagCategoryCommandCaptionGoToAddressActionSecondaryShortCuts.StringsAlt+D ShortCutL@  TAction
LockActionTagCategorySelected OperationCaption   &LåsHint   Lås markerade filer  TActionUnlockActionTagCategorySelected OperationCaption	   Lås &uppHint   Lås upp markerade filer  TAction
TipsActionTagCategoryHelpCaption
Visa &tipsHelpKeywordui_tipsHint%   Visar tips om hur du använder WinSCP
ImageIndexn  TActionChangePasswordActionTagCategorySessionCaption   Ä&ndra lösenord...HelpKeywordtask_change_passwordHint   Ändra kontolösenord  TActionPrivateKeyUploadActionTagCategorySessionCaption,&Installera den publika nyckeln i servern...HelpKeywordguide_public_keyHint;   Installera den publika nyckeln för autentisering i servern  TActionRemoteNewFileActionTagCategoryRemote Selected OperationCaption&Fil...HelpKeyword	task_editHint1   Skapa fil|Skapar ny fil och öppnas den i editorn
ImageIndexM  TAction#RemoteCalculateDirectorySizesActionTagCategoryRemote Selected OperationCaption   &Beräkna katalogstorlekarHelpKeywordui_file_panel#directory_sizesHintE   Beräkna storleken på de valda katalogerna och visa dem i filpanelenShortCut�    TActionLocalNewFileActionTagCategoryLocal Selected OperationCaption&Fil...HelpKeyword	task_editHint1   Skapa fil|Skapar ny fil och öppnas den i editorn
ImageIndexM  TActionCustomizeToolbarActionTagCategoryViewCaption   &Anpassa verktygsfältetHelpKeywordui_toolbarsHint    Visa/dölj verktygsfältsknappar  TActionRenameTabActionTagCategoryTabCaption   &Byt namn på flikenHelpKeywordui_tabs#renamingHint9   Byt namn på fliken|Ändra namnet på den aktuella fliken  TActionCurrentCopyToClipboardAction2TagCategorySelected OperationCaption&Kopiera till urklippHelpKeywordclipboard#copyHint)Kopiera de markerade filerna till urklipp
ImageIndexoShortCutC@  TActionFileColorsPreferencesActionTagCategoryViewCaption   Fil&färger...HelpKeywordui_pref_file_colorsHint   Konfigurera filfärgsregler  TAction$CurrentCopyToClipboardFocusedAction2TagCategoryFocused OperationCaption&Kopiera till urklippHelpKeywordclipboard#copyHint)Kopiera de markerade filerna till urklipp
ImageIndexoShortCutC@  TActionCommanderLocalPanelActionTagCategoryViewCaption   &Vänster panelHelpKeywordui_file_panelHint   Ändra vänster panellayout  TActionCommanderRemotePanelActionTagCategoryViewCaption   &Höger panelHelpKeywordui_file_panelHint   Ändra höger panellayout  TActionRemoteExploreDirectoryActionTagCategoryRemote DirectoryCaption&Utforska katalogHint+   Öppnar utforskaren i aktuell lokal katalog
ImageIndex8ShortCutE�    TActionLocalLocalCopyActionTag	CategoryLocal Selected OperationCaption&Kopiera...HintMKopiera den/de valda filen/filerna till en annan katalog eller ett annat namn
ImageIndexN  TActionLocalLocalMoveActionTag	CategoryLocal Selected OperationCaption
&Flytta...HintD   Flytta de valda filerna till en annan katalog eller byt namn på dem
ImageIndexd  TActionLocalOtherCopyActionTagCategoryLocal Selected OperationCaption&Kopiera...HintMKopiera den/de valda filen/filerna till en annan katalog eller ett annat namn
ImageIndexp  TActionLocalOtherMoveActionTagCategoryLocal Selected OperationCaption
&Flytta...HintD   Flytta de valda filerna till en annan katalog eller byt namn på dem
ImageIndexq  TAction"LocalCalculateDirectorySizesActionTagCategoryLocal Selected OperationCaption   &Beräkna katalogstorlekarHelpKeywordui_file_panel#directory_sizesHintE   Beräkna storleken på de valda katalogerna och visa dem i filpanelenShortCut�    TActionLocalLocalCopyFocusedActionTagCategoryLocal Focused OperationCaption&Kopiera...HintMKopiera den/de valda filen/filerna till en annan katalog eller ett annat namn
ImageIndexN  TActionLocalLocalMoveFocusedActionTagCategoryLocal Focused OperationCaption
&Flytta...HintD   Flytta de valda filerna till en annan katalog eller byt namn på dem
ImageIndexd  TActionNewTabActionTagCategoryTabCaption&Ny flikHelpKeywordui_tabs#workingHint   Öppna ny flik
ImageIndexs  TActionNewLocalTabActionTagCategoryTabCaption&Lokal flikHelpKeywordui_tabs#workingHint&   Öppna ny flik med två lokala paneler
ImageIndexsShortCutN`  TActionNewRemoteTabActionTagCategoryTabCaption   &FjärrflikHelpKeywordui_tabs#workingHint<   Öppna ny flik med en lokal panel och en fjärrsessionspanel
ImageIndexShortCutN@  TActionDefaultToNewRemoteTabActionTagCategoryTabCaption   &Standard till fjärrflikenHintc   När det är aktiverat öppnar kommandot Ny flik en ny fjärrflik. Annars öppnas en ny lokal flik.  TActionCalculateDirectorySizesActionTagCategorySelected OperationCaption   &Beräkna katalogstorlekarHelpKeywordui_file_panel#directory_sizesHintE   Beräkna storleken på de valda katalogerna och visa dem i filpanelenShortCut�    TActionLocalOtherDirActionTag	CategoryLocal DirectoryCaption   Sökväg frå&n annan panelHelpKeywordtask_navigate#special_commandsHint,   Öppna samma katalog som i den andra panelenShortCut�@  TActionRemoteOtherDirActionTagCategoryRemote DirectoryCaption   Sökväg frå&n annan panelHelpKeywordtask_navigate#special_commandsHint,   Öppna samma katalog som i den andra panelenShortCut�@  TActionIncrementalSearchStartActionTagCategoryCommandCaptionIncrementalSearchStartActionShortCutF@  TActionRemoteThumbnailActionTagCategoryStyleCaption&MiniatyrerHelpKeywordui_file_panel#view_styleHintMiniatyrer|Visa miniatyrer  TActionLocalReportActionTagCategoryStyleCaption&Detaljerad listaHelpKeywordui_file_panel#view_styleHint&Detaljerad lista|Visa detaljerad lista
ImageIndex  TActionLocalThumbnailActionTagCategoryStyleCaption&MiniatyrerHelpKeywordui_file_panel#view_styleHintMiniatyrer|Visa miniatyrer   TTBXPopupMenuExplorerBarPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left� TopP TTBXItemAddress2ActionExplorerAddressBandAction  TTBXItemStandardButtons1ActionExplorerToolbarBandAction  TTBXItemSelectionButtons1ActionExplorerSelectionBandAction  TTBXItemSessionButtons2ActionExplorerSessionBandAction2  TTBXItemPreferencesButtons1ActionExplorerPreferencesBandAction  TTBXItemSortButtons3ActionExplorerSortBandAction  TTBXItemTBXItem3ActionExplorerUpdatesBandAction  TTBXItemTBXItem4ActionExplorerTransferBandAction  TTBXItem	TBXItem16Action ExplorerCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem27  TTBXItemTBXItem7ActionLockToolbarsAction  TTBXItem	TBXItem48ActionSelectiveToolbarTextAction  TTBXSubmenuItemTBXSubmenuItem15ActionToolbarIconSizeAction TTBXItem
TBXItem127ActionToolbarIconSizeNormalAction	RadioItem	  TTBXItem
TBXItem120ActionToolbarIconSizeLargeAction	RadioItem	  TTBXItem
TBXItem128ActionToolbarIconSizeVeryLargeAction	RadioItem	   TTBXSubmenuItemTBXSubmenuItem4ActionCustomizeToolbarAction  TTBXSeparatorItemN5  TTBXItemSessionsTabs2ActionSessionsTabsAction2  TTBXItem
StatusBar2ActionStatusBarAction  TTBXSeparatorItemN72  TTBXSubmenuItemQueue7Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow6ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty6ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide5ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN71  TTBXItemToolbar5ActionQueueToolbarAction  TTBXItem	TBXItem85ActionQueueFileListAction  TTBXSeparatorItemN70  TTBXItem
Customize5ActionQueuePreferencesAction   TTBXItemTree4ActionRemoteTreeAction   TTimerSessionIdleTimerEnabledInterval�OnTimerSessionIdleTimerTimerLeft TopP  TTBXPopupMenuCommanderBarPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�Top TTBXItemCommandsButtons2ActionCommanderCommandsBandAction  TTBXItemSessionButtons5ActionCommanderSessionBandAction2  TTBXItemPreferencesButtons4ActionCommanderPreferencesBandAction  TTBXItemSortButtons2ActionCommanderSortBandAction  TTBXItemTBXItem2ActionCommanderUpdatesBandAction  TTBXItemTBXItem5ActionCommanderTransferBandAction  TTBXItem	TBXItem15Action!CommanderCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem24  TTBXItemTBXItem6ActionLockToolbarsAction  TTBXItem	TBXItem46ActionSelectiveToolbarTextAction  TTBXSubmenuItemTBXSubmenuItem14ActionToolbarIconSizeAction TTBXItem
TBXItem123ActionToolbarIconSizeNormalAction	RadioItem	  TTBXItem
TBXItem117ActionToolbarIconSizeLargeAction	RadioItem	  TTBXItem
TBXItem126ActionToolbarIconSizeVeryLargeAction	RadioItem	   TTBXSubmenuItem	TBXItem77ActionCustomizeToolbarAction  TTBXSeparatorItemN26  TTBXItemSessionsTabs1ActionSessionsTabsAction2  TTBXItemCommandLine2ActionCommandLinePanelAction  TTBXItemCommandsToolbar1ActionToolBar2Action  TTBXItem
StatusBar8ActionStatusBarAction  TTBXSeparatorItemN27  TTBXSubmenuItemLocalPanel1ActionCommanderLocalPanelAction TTBXItemHistoryButtons3Action CommanderLocalHistoryBandAction2  TTBXItemNavigationButtons3Action#CommanderLocalNavigationBandAction2  TTBXItem	TBXItem40ActionCommanderLocalFileBandAction2  TTBXItem	TBXItem43Action"CommanderLocalSelectionBandAction2  TTBXSeparatorItemN23  TTBXItemTree7ActionLocalTreeAction  TTBXSeparatorItemN77  TTBXItem
StatusBar6ActionLocalStatusBarAction2   TTBXSubmenuItemRemotePanel2ActionCommanderRemotePanelAction TTBXItemHistoryButtons4Action!CommanderRemoteHistoryBandAction2  TTBXItemNavigationButtons4Action$CommanderRemoteNavigationBandAction2  TTBXItem	TBXItem41ActionCommanderRemoteFileBandAction2  TTBXItem	TBXItem42Action#CommanderRemoteSelectionBandAction2  TTBXSeparatorItemN25  TTBXItemTree8ActionRemoteTreeAction  TTBXSeparatorItemN78  TTBXItem
StatusBar7ActionRemoteStatusBarAction2   TTBXSubmenuItemOptions1Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow5ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty5ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide4ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN69  TTBXItemToolbar4ActionQueueToolbarAction  TTBXItem	TBXItem84ActionQueueFileListAction  TTBXSeparatorItemN68  TTBXItem
Customize4ActionQueuePreferencesAction    TTBXPopupMenuRemotePanelPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left8Top TTBXSubmenuItemTBXSubmenuItem8Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem86ActionRemoteOpenDirAction  TTBXItem	TBXItem99ActionRemoteExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem13  TTBXItem	TBXItem87ActionRemoteParentDirAction  TTBXItem	TBXItem88ActionRemoteRootDirAction  TTBXItem	TBXItem89ActionRemoteHomeDirAction  TTBXItem
TBXItem109ActionRemoteOtherDirAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem90ActionRemoteBackAction  TTBXItem	TBXItem91ActionRemoteForwardAction   TTBXItem	TBXItem32ActionRemoteRefreshAction  TTBXItem	TBXItem30ActionRemoteAddBookmarkAction2  TTBXItem	TBXItem26ActionRemoteFilterAction  TTBXItemCopyPathtoClipboard1ActionRemotePathToClipboardAction2  TTBXSeparatorItemN51  TTBXItemHistoryButtons5Action!CommanderRemoteHistoryBandAction2  TTBXItemNavigationButtons5Action$CommanderRemoteNavigationBandAction2  TTBXItem	TBXItem14ActionCommanderRemoteFileBandAction2  TTBXItem	TBXItem45Action#CommanderRemoteSelectionBandAction2  TTBXSeparatorItemTBXSeparatorItem26  TTBXItem	TBXItem37ActionLockToolbarsAction  TTBXItem	TBXItem49ActionSelectiveToolbarTextAction  TTBXSubmenuItemTBXSubmenuItem13ActionToolbarIconSizeAction TTBXItem
TBXItem121ActionToolbarIconSizeNormalAction	RadioItem	  TTBXItem
TBXItem119ActionToolbarIconSizeLargeAction	RadioItem	  TTBXItem
TBXItem122ActionToolbarIconSizeVeryLargeAction	RadioItem	   TTBXSubmenuItemTBXSubmenuItem9ActionCustomizeToolbarAction  TTBXSeparatorItemN28  TTBXItemTree5ActionRemoteTreeAction  TTBXSeparatorItemN75  TTBXItem
StatusBar9ActionRemoteStatusBarAction2   TTBXPopupMenuLocalPanelPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left8TopP TTBXSubmenuItemTBXSubmenuItem10Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem92ActionLocalOpenDirAction  TTBXItem	TBXItem93ActionLocalExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem15  TTBXItem	TBXItem94ActionLocalParentDirAction  TTBXItem	TBXItem95ActionLocalRootDirAction  TTBXItem	TBXItem96ActionLocalHomeDirAction  TTBXItem
TBXItem113ActionLocalOtherDirAction  TTBXSeparatorItemTBXSeparatorItem16  TTBXItem	TBXItem97ActionLocalBackAction  TTBXItem	TBXItem98ActionLocalForwardAction   TTBXItem	TBXItem34ActionLocalRefreshAction  TTBXItem	TBXItem27ActionLocalFilterAction  TTBXItem	TBXItem31ActionLocalAddBookmarkAction2  TTBXItemCopyPathtoClipboard2ActionLocalPathToClipboardAction2  TTBXSeparatorItemN52  TTBXItemHistoryButtons6Action CommanderLocalHistoryBandAction2  TTBXItemNavigationButtons6Action#CommanderLocalNavigationBandAction2  TTBXItem	TBXItem39ActionCommanderLocalFileBandAction2  TTBXItem	TBXItem44Action"CommanderLocalSelectionBandAction2  TTBXSeparatorItemTBXSeparatorItem25  TTBXItem	TBXItem38ActionLockToolbarsAction  TTBXItem	TBXItem47ActionSelectiveToolbarTextAction  TTBXSubmenuItemTBXSubmenuItem16ActionToolbarIconSizeAction TTBXItem
TBXItem129ActionToolbarIconSizeNormalAction	RadioItem	  TTBXItem
TBXItem118ActionToolbarIconSizeLargeAction	RadioItem	  TTBXItem
TBXItem130ActionToolbarIconSizeVeryLargeAction	RadioItem	   TTBXSubmenuItemTBXSubmenuItem6ActionCustomizeToolbarAction  TTBXSeparatorItemN29  TTBXItemTree6ActionLocalTreeAction  TTBXSeparatorItemN76  TTBXItemStatusBar10ActionLocalStatusBarAction2   TTBXPopupMenuLocalDirViewColumnPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left� TopX TTBXItemSortAscending1ActionSortColumnAscendingAction  TTBXItemSortDescending1ActionSortColumnDescendingAction  TTBXItemLocalSortByExtColumnPopupItemActionLocalSortByExtAction2  TTBXItemHidecolumn1ActionHideColumnAction  TTBXSeparatorItemN37  TTBXSubmenuItemLocalFormatSizeBytesPopupItemCaptionVisa &filstorlekar iHelpKeywordui_pref_panels#commonHint$   Välj visningsformat för filstorlek TTBXItem	TBXItem64ActionFormatSizeBytesNoneAction  TTBXItem	TBXItem65ActionFormatSizeBytesKilobytesAction  TTBXItem	TBXItem66ActionFormatSizeBytesShortAction   TTBXItem%LocalCalculateDirectorySizesPopupItemAction"LocalCalculateDirectorySizesAction  TTBXSeparatorItemTBXSeparatorItem8  TTBXSubmenuItemLocalColumnsSubmenuItemCaption	&KolumnerHelpKeywordui_file_panel#selecting_columns TTBXItemName3ActionShowHideLocalNameColumnAction2  TTBXItemSize3ActionShowHideLocalSizeColumnAction2  TTBXItemType2ActionShowHideLocalTypeColumnAction2  TTBXItemModification3Action!ShowHideLocalChangedColumnAction2  TTBXItemAttributes3ActionShowHideLocalAttrColumnAction2  TTBXSeparatorItemTBXSeparatorItem73  TTBXItem
TBXItem264ActionAutoSizeLocalColumnsAction  TTBXItem
TBXItem112ActionResetLayoutLocalColumnsAction    TTBXPopupMenuRemoteDirViewColumnPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�TopX TTBXItem	MenuItem1ActionSortColumnAscendingAction	RadioItem	  TTBXItem	MenuItem2ActionSortColumnDescendingAction	RadioItem	  TTBXItemRemoteSortByExtColumnPopupItemActionRemoteSortByExtAction2  TTBXItemHidecolumn2ActionHideColumnAction  TTBXSeparatorItemN38  TTBXSubmenuItemRemoteFormatSizeBytesPopupItemCaptionVisa &filstorlekar iHelpKeywordui_pref_panels#commonHint$   Välj visningsformat för filstorlek TTBXItem	TBXItem67ActionFormatSizeBytesNoneAction  TTBXItem	TBXItem53ActionFormatSizeBytesKilobytesAction  TTBXItem	TBXItem55ActionFormatSizeBytesShortAction   TTBXItem&RemoteCalculateDirectorySizesPopupItemAction#RemoteCalculateDirectorySizesAction  TTBXSeparatorItemTBXSeparatorItem7  TTBXSubmenuItemRemoteColumnsSubmenuItemCaption	&KolumnerHelpKeywordui_file_panel#selecting_columns TTBXItemName4ActionShowHideRemoteNameColumnAction2  TTBXItemSize4ActionShowHideRemoteSizeColumnAction2  TTBXItemTBXItem8ActionShowHideRemoteTypeColumnAction2  TTBXItemModification4Action"ShowHideRemoteChangedColumnAction2  TTBXItemPermissions1Action!ShowHideRemoteRightsColumnAction2  TTBXItemOwner2Action ShowHideRemoteOwnerColumnAction2  TTBXItemGroup2Action ShowHideRemoteGroupColumnAction2  TTBXItemTBXItem1Action%ShowHideRemoteLinkTargetColumnAction2  TTBXSeparatorItemTBXSeparatorItem20  TTBXItem
TBXItem114ActionAutoSizeRemoteColumnsAction  TTBXItem
TBXItem115ActionResetLayoutRemoteColumnsAction    TTBXPopupMenu
QueuePopupImagesGlyphsModule.ExplorerImagesOnPopupQueuePopupPopupOptionstboShowHint LefthTop�  TTBXItem
ShowQuery1ActionQueueItemQueryAction  TTBXItem
ShowError1ActionQueueItemErrorAction  TTBXItemShowPrompt1ActionQueueItemPromptAction  TTBXSeparatorItemN53  TTBXItemExecuteNow1ActionQueueItemExecuteAction  TTBXItemTBXItem9ActionQueueItemPauseAction  TTBXItem	TBXItem10ActionQueueItemResumeAction  TTBXItemDelete4ActionQueueItemDeleteAction  TTBXComboBoxItemQueuePopupSpeedComboBoxItemActionQueueItemSpeedAction	ShowImage	OnAdjustImageIndex+QueuePopupSpeedComboBoxItemAdjustImageIndex  TTBXSeparatorItemN54  TTBXItemMoveUp1ActionQueueItemUpAction  TTBXItem	MoveDown1ActionQueueItemDownAction  TTBXSeparatorItemN67  TTBXItemQueueEnableItemActionQueueEnableAction  TTBXSubmenuItemTBXSubmenuItem1Caption&AllaHelpKeywordui_queue#manageHint&   Administrationskommandon för kömassa TTBXItem	TBXItem11ActionQueuePauseAllAction  TTBXItem	TBXItem12ActionQueueResumeAllAction  TTBXItem
TBXItem142ActionQueueDeleteAllAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem51ActionQueueDeleteAllDoneAction   TTBXSubmenuItemTBXSubmenuItem3ActionQueueCycleOnceEmptyActionDropdownCombo	 TTBXItem	TBXItem28ActionQueueIdleOnceEmptyAction	RadioItem	  TTBXItem	TBXItem13ActionQueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem	TBXItem68ActionQueueSuspendOnceEmptyAction2	RadioItem	  TTBXItem	TBXItem29ActionQueueShutDownOnceEmptyAction2	RadioItem	   TTBXSubmenuItemQueue2Caption&AlternativHelpKeywordui_queueHint   Konfigurera kölista TTBXItemShow4ActionQueueShowAction	RadioItem	  TTBXItemHidewhenEmpty4ActionQueueHideWhenEmptyAction	RadioItem	  TTBXItemHide3ActionQueueHideAction	RadioItem	  TTBXSeparatorItemN66  TTBXItemToolbar3ActionQueueToolbarAction  TTBXItem	TBXItem83ActionQueueFileListAction  TTBXSeparatorItemTBXSeparatorItem23  TTBXItem
TBXItem116ActionQueueResetLayoutColumnsAction  TTBXSeparatorItemN65  TTBXItem
Customize3ActionQueuePreferencesAction    TTBXPopupMenuRemoteDirViewPopup	AutoPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint LefthTop� TTBXSubmenuItemGoTo4Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemOpenDirectoryBookmark3ActionRemoteOpenDirAction  TTBXItem
TBXItem100ActionRemoteExploreDirectoryAction  TTBXSeparatorItemN81  TTBXItemParentDirectory4ActionRemoteParentDirAction  TTBXItemRootDirectory4ActionRemoteRootDirAction  TTBXItemHomeDirectory4ActionRemoteHomeDirAction  TTBXSeparatorItemN80  TTBXItemBack4ActionRemoteBackAction  TTBXItemForward4ActionRemoteForwardAction   TTBXItemRefresh4ActionRemoteRefreshAction  TTBXItemAddToBookmarks4ActionRemoteAddBookmarkAction2  TTBXItem	TBXItem35ActionRemoteFilterAction  TTBXItemCopyPathtoClipboard6ActionRemotePathToClipboardAction2  TTBXSeparatorItemN79  TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135ActionNewFileAction  TTBXItem
TBXItem136ActionNewDirAction  TTBXItem
TBXItem209ActionNewLinkAction   TTBXItem	TBXItem75ActionPasteAction3  TTBXSubmenuItem$RemoteDirViewPopupCustomCommandsMenuActionCustomCommandsNonFileAction   TTBXPopupMenuLocalDirViewPopup	AutoPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�Top� TTBXSubmenuItemGoTo5Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemOpenDirectoryBookmark4ActionLocalOpenDirAction  TTBXItemExploreDirectory2ActionLocalExploreDirectoryAction  TTBXSeparatorItemN84  TTBXItemParentDirectory5ActionLocalParentDirAction  TTBXItemRootDirectory5ActionLocalRootDirAction  TTBXItemHomeDirectory5ActionLocalHomeDirAction  TTBXSeparatorItemN83  TTBXItemBack5ActionLocalBackAction  TTBXItemForward5ActionLocalForwardAction   TTBXItemRefresh5ActionLocalRefreshAction  TTBXItem	TBXItem36ActionLocalFilterAction  TTBXItemAddToBookmarks5ActionLocalAddBookmarkAction2  TTBXItemCopyPathtoClipboard7ActionLocalPathToClipboardAction2  TTBXSeparatorItemN82  TTBXSubmenuItemTBXSubmenuItem7Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem	TBXItem70ActionNewFileAction  TTBXItem	TBXItem71ActionNewDirAction   TTBXItem	TBXItem76ActionPasteAction3   TTBXPopupMenuRemoteAddressPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left� Top� TTBXItem	TBXItem33ActionRemoteRefreshAction  TTBXItem	TBXItem24ActionRemoteAddBookmarkAction2  TTBXItem	TBXItem25ActionRemotePathToClipboardAction2  TTBXSeparatorItemTBXSeparatorItem1  TTBXItem	TBXItem17ActionRemoteOpenDirAction  TTBXSubmenuItemTBXSubmenuItem2Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem18ActionRemoteParentDirAction  TTBXItem	TBXItem19ActionRemoteRootDirAction  TTBXItem	TBXItem20ActionRemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItem	TBXItem21ActionRemoteBackAction  TTBXItem	TBXItem22ActionRemoteForwardAction    TTBXPopupMenuSessionsPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left�Top�  TTBXItem
TBXItem124ActionCloseTabAction  TTBXItem
TBXItem219ActionDuplicateTabAction  TTBXItem	TBXItem78ActionRenameTabAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXColorItemColorMenuItemActionColorMenuAction2ColorclNone  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem	TBXItem79ActionDisconnectSessionAction  TTBXItem	TBXItem80ActionReconnectSessionAction  TTBXItem
TBXItem125ActionSaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem56ActionFileSystemInfoAction  TTBXItem	TBXItem52ActionSessionGenerateUrlAction2  TTBXSeparatorItemTBXSeparatorItem34  TTBXSubmenuItemSessionsNewTabItemActionNewTabActionDropdownCombo	 TTBXItem
TBXItem104ActionNewRemoteTabAction  TTBXItem
TBXItem105ActionNewLocalTabAction  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem
TBXItem106ActionDefaultToNewRemoteTabAction   TTBXSubmenuItemTBXSubmenuItem23ActionSavedSessionsAction2OptionstboDropdownArrow   TTBXSeparatorItemTBXSeparatorItem35  TTBXItemSessionsTabs4ActionSessionsTabsAction2   TTBXPopupMenuLocalFilePopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint LeftTopP TTBXItemLocalOpenMenuItemActionCurrentOpenAction  TTBXSubmenuItemLocalEditMenuItemActionCurrentEditFocusedActionDropdownCombo	OnPopupFocusedEditMenuItemPopup  TTBXSubmenuItemLocalCopyMenuItemActionLocalCopyFocusedActionDropdownCombo	 TTBXItem	TBXItem73ActionLocalCopyFocusedNonQueueAction  TTBXItem	TBXItem74ActionLocalCopyFocusedQueueAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem54ActionLocalMoveFocusedAction   TTBXItemLocalLocalCopyMenuItemActionLocalLocalCopyFocusedAction  TTBXItem
TBXItem101ActionLocalLocalMoveFocusedAction  TTBXItem	TBXItem57ActionCurrentDeleteFocusedAction  TTBXItem	TBXItem58ActionCurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem81Action$CurrentCopyToClipboardFocusedAction2  TTBXSeparatorItemTBXSeparatorItem3  TTBXSubmenuItem LocalFilePopupCustomCommandsMenuActionCustomCommandsFileAction TTBXItem    TTBXSubmenuItemTBXSubmenuItem5Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem59ActionFileListToCommandLineAction  TTBXItem	TBXItem60ActionFileListToClipboardAction  TTBXItem	TBXItem61ActionFullFileListToClipboardAction   TTBXSeparatorItemTBXSeparatorItem4  TTBXItem	TBXItem63ActionCurrentPropertiesFocusedAction  TTBXItem	TBXItem50ActionCurrentSystemMenuFocusedAction   TTBXPopupMenuLocalBrowserPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left(Top�  TTBXItem	TBXItem62ActionCloseTabAction  TTBXItem
TBXItem102ActionDuplicateTabAction  TTBXItem
TBXItem103ActionRenameTabAction  TTBXSeparatorItemTBXSeparatorItem21  TTBXSubmenuItemTBXSubmenuItem12ActionNewTabActionDropdownCombo	 TTBXItem
TBXItem107ActionNewRemoteTabAction  TTBXItem
TBXItem108ActionNewLocalTabAction  TTBXSeparatorItemTBXSeparatorItem19  TTBXItem
TBXItem111ActionDefaultToNewRemoteTabAction   TTBXSubmenuItemTBXSubmenuItem11ActionSavedSessionsAction2OptionstboDropdownArrow   TTBXSeparatorItemTBXSeparatorItem22  TTBXItem
TBXItem110ActionSessionsTabsAction2   TTBXPopupMenuNewTabPopupImagesGlyphsModule.ExplorerImagesOptionstboShowHint Left Top�  TTBXItemNewRemoteTabItemActionNewRemoteTabAction  TTBXItemNewLocalTabItemActionNewLocalTabAction  TTBXSeparatorItemTBXSeparatorItem67  TTBXItem
TBXItem232ActionDefaultToNewRemoteTabAction     TPF0TOpenDirectoryDialogOpenDirectoryDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_opendirBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionOpen directoryClientHeightVClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnShowFormShow
DesignSize�V 
TextHeight TLabel	EditLabelLeft.TopWidthRHeightCaption   &Öppna katalog:  TImageImageLeftTopWidth Height AutoSize	  THistoryComboBoxLocalDirectoryEditLeft.TopWidth6HeightAnchorsakLeftakTopakRight TabOrderTextLocalDirectoryEditOnChangeDirectoryEditChangeSaveOn   THistoryComboBoxRemoteDirectoryEditLeft.TopWidth�HeightAnchorsakLeftakTopakRight DropDownCount	MaxLength�TabOrder TextRemoteDirectoryEditOnChangeDirectoryEditChangeSaveOn   TButtonOKBtnLeft� Top5WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeftTop5WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeftTop7Width�Height� 
ActivePageSessionBookmarksSheetAnchorsakLeftakTopakRightakBottom TabOrderOnChangePageControlChange 	TTabSheetSessionBookmarksSheetTagCaption   Sessionsbokmärken
DesignSize��   TListBoxSessionBookmarksListTagLeftTopWidthHHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSessionBookmarkButtonTagLeftSTopWidthPHeightAnchorsakTopakRight Caption   &Lägg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSessionBookmarkButtonTagLeftSTop$WidthPHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSessionBookmarkButtonTag�LeftSTop� WidthPHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSessionBookmarkButtonTagLeftSTop� WidthPHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick   	TTabSheetSharedBookmarksSheetTagCaption   Delade bokmärken
ImageIndex
DesignSize��   TListBoxSharedBookmarksListTagLeftTopWidthHHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClickBookmarksListClick
OnDblClickBookmarksListDblClick
OnDragDropBookmarksListDragDrop
OnDragOverBookmarksListDragOver	OnEndDragBookmarksListEndDrag	OnKeyDownBookmarksListKeyDownOnStartDragBookmarksListStartDrag  TButtonAddSharedBookmarkButtonTagLeftSTopWidthPHeightAnchorsakTopakRight Caption   &Lägg tillTabOrderOnClickAddBookmarkButtonClick  TButtonRemoveSharedBookmarkButtonTagLeftSTop$WidthPHeightAnchorsakTopakRight Caption&Ta bortTabOrderOnClickRemoveBookmarkButtonClick  TButtonUpSharedBookmarkButtonTag�LeftSTop� WidthPHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickBookmarkButtonClick  TButtonDownSharedBookmarkButtonTagLeftSTop� WidthPHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickBookmarkButtonClick  TButtonShortCutSharedBookmarkButtonTagLeftSTopCWidthPHeightAnchorsakTopakRight Caption   &Genväg...TabOrderOnClickShortCutBookmarkButtonClick    TButtonLocalDirectoryBrowseButtonLeftjTopWidthPHeightAnchorsakTopakRight Caption   Blädd&ra...TabOrderOnClickLocalDirectoryBrowseButtonClick  TButtonSwitchButtonLeftTop5Width� HeightAnchorsakLeftakBottom CaptionP&latsprofiler...ModalResultTabOrderOnClickSwitchButtonClick  TButton
HelpButtonLeftjTop5WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick      TPF0TPreferencesDialogPreferencesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_preferencesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption   InställningarClientHeight9ClientWidth]Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnCloseQueryFormCloseQuery
OnShortCutFormShortCutOnShowFormShow
DesignSize]9 
TextHeight TButtonOKButtonLeftYTop�WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCloseButtonLeft�Top�WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPanel	MainPanelLeft Top Width]Height�AlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  TPageControlPageControlLeft� Top Width�Height�
ActivePagePreferencesSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheetPreferencesSheetTagHelpType	htKeywordHelpKeywordui_pref_environmentCaption   Miljö
ImageIndex
TabVisible
DesignSize��  	TGroupBoxCommonPreferencesGroupLeftTopWidth�Height0AnchorsakLeftakTopakRight Caption   BekräftelserTabOrder 
DesignSize�0  	TCheckBoxSynchronizeSummaryCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption   &SynkroniseringsöversiktTabOrder
OnClickControlChange  	TCheckBoxConfirmOverwritingCheckLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption   Ö&verskrivning av filerTabOrderOnClickControlChange  	TCheckBoxConfirmDeletingCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption%&Borttagning av filer (rekommenderad)TabOrderOnClickControlChange  	TCheckBoxConfirmClosingSessionCheck2LeftTop� Width�HeightAnchorsakLeftakTopakRight Caption*   Stäng sessioner när programmet avs&lutasTabOrderOnClickControlChange  	TCheckBoxDDTransferConfirmationCheck2LeftTop-Width�HeightAnchorsakLeftakTopakRight Caption?   D&ra && släpp operationer och klistra in i andra applikationerTabOrderOnClickControlChange  	TCheckBoxContinueOnErrorCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption*   Fortsätt vid &fel (avancerade användare)TabOrderOnClickControlChange  	TCheckBoxConfirmExitOnCompletionCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption.   Avsluta a&pplikationen vid slutförd operationTabOrderOnClickControlChange  	TCheckBoxConfirmResumeCheckLeftTop[Width�HeightAnchorsakLeftakTopakRight Caption   &Återuppta överföringTabOrderOnClickControlChange  	TCheckBoxConfirmCommandSessionCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption   Öppna separat &skalsessionTabOrder	OnClickControlChange  	TCheckBoxConfirmRecyclingCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption &Flytta filer till papperskorgenTabOrderOnClickControlChange  	TCheckBoxConfirmTransferringCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   &Överföring av filerTabOrder OnClickControlChange  TStaticTextBackgroundConfirmationsLinkLeftToprWidth�Height	AlignmenttaRightJustifyAnchorsakLeftakTopakRight AutoSizeCaption/   Ändra bekräftelser av bakgrundsöverföringarTabOrderTabStop	OnClick BackgroundConfirmationsLinkClick   	TGroupBoxNotificationsGroupLeftTop8Width�HeightHAnchorsakLeftakTopakRight CaptionMeddelandenTabOrder
DesignSize�H  TLabelBeepOnFinishAfterTextLeft�TopWidthHeightAnchorsakTopakRight CaptionsShowAccelChar  	TCheckBoxBeepOnFinishCheckLeftTopWidthMHeightAnchorsakLeftakTopakRight Caption=   S&ystemljud när operationen är klar, om den pågår mer änTabOrder OnClickControlChange  TUpDownEditBeepOnFinishAfterEditLeft^TopWidthIHeight	AlignmenttaRightJustify	Increment       �@MaxValue      ��@AnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChange  	TCheckBoxBalloonNotificationsCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight CaptionK   Visa ballong&meddelanden i aktivitetsfältets statusområde (systemfältet)TabOrderOnClickControlChange    	TTabSheetLogSheetTagHelpType	htKeywordHelpKeywordui_pref_loggingCaptionLoggning
ImageIndex
TabVisible
DesignSize��  TLabelLogProtocolHintLabelLeftTop+Width�Height+AnchorsakLeftakTopakRight AutoSizeCaption^   Den valda loggningsnivån försämrar prestandan kraftigt. Använd den endast vid felsökning.ShowAccelCharWordWrap	  	TGroupBoxLoggingGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Alternativ för loggningTabOrder 
DesignSize��   TLabelLogMaxSizeCountFilesLabelLeftTop� WidthHeightAnchorsakTopakRight CaptionfilerFocusControlLogMaxSizeCountEditShowAccelChar  TLabelLogFileNameLabelLeftTop-Width2HeightCaption   &Loggsökväg:FocusControlLogFileNameEdit3OnClickControlChange  TFilenameEditLogFileNameEdit3LeftTop?Width�HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogKinddkSave
DefaultExtlogFilter4Sessionsloggfilar (*.log)|*.log|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för sessionslogg.ClickKey@AnchorsakLeftakTopakRight TabOrderTextLogFileNameEdit3OnChangeControlChange  TPanelLogFilePanelLeftTopVWidthAHeightAnchorsakLeftakTopakRight 
BevelOuterbvNoneTabOrder TRadioButtonLogFileAppendButtonLeft TopWidthtHeightCaption   L&ägg tillTabOrder OnClickControlChange  TRadioButtonLogFileOverwriteButtonLeftzTopWidthtHeightCaption   Sk&riv överTabOrderOnClickControlChange   	TComboBoxLogProtocolCombo2Left1TopWidth� HeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChangeControlChangeItems.Strings	ReduceradNormalDebug 1Debug 2   TStaticTextLogFileNameHintTextLeft1TopTWidth� Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  	TCheckBoxEnableLoggingCheckLeftTopWidth HeightAnchorsakLeftakTopakRight Caption!   Aktivera &sessionslogg på nivå:TabOrder OnClickControlChange  	TCheckBoxLogSensitiveCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption/   Logga &lösenord och annan känslig informationTabOrder	OnClickControlChange  	TCheckBoxLogMaxSizeCheckLeftTopqWidthHeightAnchorsakLeftakTopakRight Caption$   &Rotera loggfiler efter de har nåttTabOrderOnClickControlChange  	TComboBoxLogMaxSizeComboLeft1TopnWidth� HeightAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeOnExitSizeComboExitItems.Strings1M10M100M1G   	TCheckBoxLogMaxSizeCountCheckLeft-Top� Width� HeightAnchorsakLeftakTopakRight Caption!   &Ta bort gamla loggfiler, behållTabOrderOnClickControlChange  TUpDownEditLogMaxSizeCountEditLeft1Top� WidthHHeightMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrderOnChangeControlChange   	TGroupBoxActionsLoggingGroupLeftTop� Width�HeightZAnchorsakLeftakTopakRight CaptionXML-loggTabOrder
DesignSize�Z  TFilenameEditActionsLogFileNameEditLeftTop-Width�HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogKinddkSave
DefaultExtxmlFilter0XML-loggfiler (*.xml)|*.xml|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för XML-logg.ClickKey@AnchorsakLeftakTopakRight TabOrderTextActionsLogFileNameEditOnChangeControlChange  TStaticTextActionsLogFileNameHintTextLeft1TopBWidth� Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   möns&terTabOrderTabStop	  	TCheckBoxEnableActionsLoggingCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionAktivera &XML-logg till fil:TabOrder OnClickControlChange    	TTabSheetGeneralSheetTagHelpType	htKeywordHelpKeywordui_pref_interfaceCaption   Gränssnitt
ImageIndex
TabVisible
DesignSize��  TLabelInterfaceChangeLabelLeftTopWidth� HeightCaption.   Ändringar kommer att gälla vid nästa start.ShowAccelChar  	TGroupBoxInterfaceGroupLeftTop<Width�Height� AnchorsakLeftakTopakRight Caption   AnvändargränssnittTabOrder
DesignSize��   TLabelCommanderDescriptionLabel2Left� TopWidth!HeightsAnchorsakLeftakTopakRight AutoSizeCaption�   - två paneler (vänster för lokal katalog, höger för fjärrkatalog)
- snabbkommandon som i Norton Commander (och andra liknande program som Total Commander, Midnight Commander...)
- dra && släpp till/från båda panelernaFocusControlCommanderInterfaceButton2WordWrap	OnClickCommanderClick  TLabelExplorerDescriptionLabelLeft� Top� Width!HeightCAnchorsakLeftakTopakRight AutoSizeCaptionK   - endast fjärrkatalog
- snabbkommandon som i Utforskaren
- dra && släppFocusControlExplorerInterfaceButton2WordWrap	OnClickExplorerClick  TImageCommanderInterfacePictureLeft7Top-Width Height AutoSize	OnClickCommanderClick  TImageExplorerInterfacePictureLeft7Top� Width Height AutoSize	OnClickExplorerClick  TRadioButtonCommanderInterfaceButton2LeftTopWidthtHeightCaption
&CommanderChecked	TabOrder TabStop	OnClickControlChange  TRadioButtonExplorerInterfaceButton2LeftTop� WidthoHeightCaption&UtforskareTabOrderOnClickControlChange   	TGroupBox
ThemeGroupLeftTopWidth�Height4AnchorsakLeftakTopakRight CaptionTemaTabOrder 
DesignSize�4  TLabelLabel7Left	TopWidthVHeightCaption   Gränssnitts&tema:FocusControl
ThemeCombo  	TComboBox
ThemeComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder Items.Strings
AutomatiskLjus   Mörk     	TTabSheetPanelsSheetTagHelpType	htKeywordHelpKeywordui_pref_panelsCaptionPaneler
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPanelsCommonGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   AllmäntTabOrder 
DesignSize��   TLabelLabel1Left	Top� Width[HeightCaptionVisa &filstorlek i:FocusControlFormatSizeBytesComboOnClickControlChange  TLabelLabel2Left	Top� WidthgHeightCaption   &Inkrementell sökning:FocusControlPanelSearchComboOnClickControlChange  	TCheckBoxShowHiddenFilesCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionVi&sa dolda filer (CTRL+ALT+H)TabOrder OnClickControlChange  	TCheckBoxDefaultDirIsHomeCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption!   Standardkatalog är &hemkatalogenTabOrderOnClickControlChange  	TCheckBoxPreservePanelStateCheckLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption4   Kom i&håg panelens' tillstånd när session växlasTabOrderOnClickControlChange  	TCheckBoxRenameWholeNameCheckLeftTop[Width�HeightAnchorsakLeftakTopakRight Caption&   Välj &hela namnet när filen döps omTabOrderOnClickControlChange  	TCheckBoxFullRowSelectCheckLeftToprWidth�HeightAnchorsakLeftakTopakRight Caption   Välja med h&ela radenTabOrderOnClickControlChange  	TComboBoxFormatSizeBytesComboLeft<Top� WidthxHeightStylecsDropDownListAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeItems.StringsByteKilobyteKort format   	TCheckBox!NaturalOrderNumericalSortingCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption0   Använd &numerisk sortering med naturlig ordningTabOrderOnClickControlChange  	TComboBoxPanelSearchComboLeft� Top� Width� HeightStylecsDropDownListAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeItems.Strings   Endast början av namnetAlla delar av namnetAlla kolumner   	TCheckBox AlwaysSortDirectoriesByNameCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption$Sortera alltid &kataloger efter namnTabOrderOnClickControlChange   	TGroupBoxDoubleClickGroupLeftTop� Width�HeightKAnchorsakLeftakTopakRight CaptionDubbelklickTabOrder
DesignSize�K  TLabelDoubleClickActionLabelLeft	TopWidth� HeightAnchorsakLeftakTopakRight Caption'   &Operation att utföra vid dubbelklick:FocusControlDoubleClickActionCombo  	TCheckBox"CopyOnDoubleClickConfirmationCheckLeftTop0Width�HeightAnchorsakLeftakTopakRight Caption,   &Bekräfta kopiera vid dubbelklicksoperationTabOrderOnClickControlChange  	TComboBoxDoubleClickActionComboLeft<TopWidthxHeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChangeControlChangeItems.Strings   ÖppnaKopieraRedigera    	TGroupBoxPanelFontGroupLeftTopNWidth�HeightPAnchorsakLeftakTopakRight CaptionPanel teckensnittTabOrder
DesignSize�P  TLabelPanelFontLabelLeft� TopWidthHeight0AnchorsakLeftakTopakRightakBottom AutoSizeCaptionPanelFontLabelColorclWindowParentColorShowAccelCharTransparentWordWrap	
OnDblClickPanelFontLabelDblClick  TButtonPanelFontButtonLeft	Top-Width� HeightCaption   Välj tecke&nsnittTabOrderOnClickPanelFontButtonClick  	TCheckBoxPanelFontCheckLeftTopWidth� HeightCaption   Använd anpassad &teckensnittTabOrder OnClickControlChange    	TTabSheetCommanderSheetTagHelpType	htKeywordHelpKeywordui_pref_commanderCaption	Commander
ImageIndex
TabVisible
DesignSize��  TLabelLabel3LeftTopWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaptionV   Inställningar på den här fliken gäller endast för Norton Commander-gränssnittet.ShowAccelCharWordWrap	  	TGroupBoxPanelsGroupLeftTop"Width�HeightcAnchorsakLeftakTopakRight CaptionPanelerTabOrder 
DesignSize�c  TLabelLabel8Left	TopWidth|HeightCaptionVal av &utforskarstil:FocusControlNortonLikeModeCombo  	TCheckBoxSwappedPanelsCheckLeftTop0Width�HeightAnchorsakLeftakTopakRight Caption6   B&yt paneler (lokal till höger, fjärr till vänster)TabOrderOnClickControlChange  	TComboBoxNortonLikeModeComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeItems.StringsAldrigBara musMus och tangentbord   	TCheckBoxTreeOnLeftCheckLeftTopGWidth�HeightAnchorsakLeftakTopakRight Caption(   Visa &katalogträd vänster om fillistanTabOrderOnClickControlChange   	TGroupBoxCommanderMiscGroupLeftTop� Width�HeightKAnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize�K  TLabelLabel10Left	TopWidthfHeightCaption&KortkommandonFocusControlExplorerKeyboardShortcutsCombo  	TCheckBoxUseLocationProfilesCheckLeftTop0Width�HeightAnchorsakLeftakTopakRight Caption7   &Använd platsprofiler istället för katalogbokmärkenTabOrderOnClickControlChange  	TComboBoxExplorerKeyboardShortcutsComboLeft� TopWidth� HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeItems.Strings	CommanderUtforskaren    	TGroupBoxCompareCriterionsGroupLeftTop� Width�HeightHAnchorsakLeftakTopakRight Caption   Jämför katalogkriteriumTabOrder
DesignSize�H  	TCheckBoxCompareByTimeCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Jämför efter &tidTabOrder OnClickControlChange  	TCheckBoxCompareBySizeCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption   Jämför efter &storlekTabOrderOnClickControlChange    	TTabSheetExplorerSheetTagHelpType	htKeywordHelpKeywordui_pref_explorerCaptionUtforskaren
ImageIndex
TabVisible
DesignSize��  TLabelLabel4LeftTopWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaptionM   Inställningar på den här fliken gäller endast för utforskargränssnittetShowAccelCharWordWrap	  	TGroupBox	GroupBox2LeftTop"Width�Height1AnchorsakLeftakTopakRight CaptionVisaTabOrder 
DesignSize�1  	TCheckBoxShowFullAddressCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption2   Vi&sa den fullständiga sökvägen i adressfältetTabOrder OnClickControlChange    	TTabSheetEditorSheetTagHelpType	htKeywordHelpKeywordui_pref_editorCaptionEditor
ImageIndex
TabVisible
DesignSize��  	TGroupBoxEditorPreferenceGroupLeftTopWidth�Height�AnchorsakLeftakTopakRightakBottom Caption   EditorinställningarTabOrder 
DesignSize��  	TListViewEditorListView3Left	TopWidth�HeightBAnchorsakLeftakTopakRightakBottom ColumnsCaptionEditorWidth�  CaptionMaskWidthF CaptionTextWidth-  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder 	ViewStylevsReportOnDataEditorListView3Data
OnDblClickEditorListView3DblClick	OnEndDragListViewEndDrag
OnDragDropEditorListView3DragDrop
OnDragOverListViewDragOver	OnKeyDownEditorListView3KeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddEditorButtonLeft	Top^WidthZHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddEditEditorButtonClick  TButtonEditEditorButtonLeftiTop^WidthZHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickAddEditEditorButtonClick  TButtonUpEditorButtonLeftZTop^WidthZHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownEditorButtonClick  TButtonDownEditorButtonLeftZTop}WidthZHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownEditorButtonClick  TButtonRemoveEditorButtonLeft	Top}WidthZHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveEditorButtonClick   	TGroupBoxEditingOptionsGroupLeftTop�Width�Height1AnchorsakLeftakRightakBottom CaptionRedigeringsalternativTabOrder
DesignSize�1  	TCheckBoxEditorCheckNotModifiedCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionQ   &Kontrollera att den redigerade fjärrfilen inte har ändrats innan du sparar denTabOrder OnClickControlChange    	TTabSheetIntegrationSheetTag	HelpType	htKeywordHelpKeywordui_pref_integrationCaptionIntegrering
ImageIndex
TabVisible
DesignSize��  	TGroupBoxShellIconsGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionWindowsskalTabOrder 
DesignSize��   TButtonDesktopIconButtonLeft	TopWidth�HeightAnchorsakLeftakTopakRight Caption   Skapa en ikon på skrivbor&detTabOrder OnClickIconButtonClick  TButtonSendToHookButtonLeft	Top5Width�HeightAnchorsakLeftakTopakRight CaptionB   Skapa genväg för överföring i utforskarens '&Skicka till'-menyTabOrderOnClickIconButtonClick  TButtonRegisterAsUrlHandlersButtonLeft	TophWidth�HeightAnchorsakLeftakTopakRight Caption)   Registrera för att hantera &URL-adresserTabOrderOnClick RegisterAsUrlHandlersButtonClick  TButtonAddSearchPathButtonLeft	Top� Width�HeightAnchorsakLeftakTopakRight Caption7   Lägg till sökvägen till WinSCP i miljövaribeln PATHTabOrderOnClickAddSearchPathButtonClick  TStaticTextShellIconsText2LeftjTopQWidthJHeightHint   För att lägga till genvägar, som direkt öppnar webbplats, använd ikonkommandon i 'Hantera'-menyn i dialogrutan inloggning.	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaptionAssociera ikoner med webbplatsTabOrderTabStop	    	TTabSheetCustomCommandsSheetTag
HelpType	htKeywordHelpKeywordui_pref_commandsCaption	Kommandon
ImageIndex	
TabVisible
DesignSize��  	TGroupBoxCustomCommandsGroupLeftTopWidth�Height�AnchorsakLeftakTopakRightakBottom CaptionEgna kommandonTabOrder 
DesignSize��  	TListViewCustomCommandsViewLeft	TopWidth�HeightyAnchorsakLeftakTopakRightakBottom ColumnsCaptionBeskrivningWidthU CaptionKommandoWidth�  CaptionL/FWidth#  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedParentShowHintShowHint	TabOrder 	ViewStylevsReportOnDataCustomCommandsViewData
OnDblClickCustomCommandsViewDblClick	OnEndDragListViewEndDrag
OnDragDropCustomCommandsViewDragDrop
OnDragOverCustomCommandsViewDragOver	OnKeyDownCustomCommandsViewKeyDownOnMouseMoveCustomCommandsViewMouseMoveOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCommandButtonLeft	Top�WidthdHeightAnchorsakLeftakBottom Caption   &Lägg till...StylebsSplitButtonTabOrderOnClickAddCommandButtonClickOnDropDownClickAddCommandButtonDropDownClick  TButtonRemoveCommandButtonLeft	Top�WidthdHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveCommandButtonClick  TButtonUpCommandButtonLeftZTop�WidthZHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCommandButtonClick  TButtonDownCommandButtonLeftZTop�WidthZHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCommandButtonClick  TButtonEditCommandButtonLeftsTop�WidthdHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickEditCommandButtonClick  TButtonConfigureCommandButtonLeftsTop�WidthdHeightAnchorsakLeftakBottom Caption&Konfigurera...TabOrderOnClickConfigureCommandButtonClick    	TTabSheetDragDropSheetTagHelpType	htKeywordHelpKeywordui_pref_dragdropCaption   Dra & släpp
ImageIndex

TabVisible
DesignSize��  	TGroupBoxDragDropDownloadsGroupLeftTopWidth�HeightIAnchorsakLeftakTopakRight Caption   Dra && släpp nerladdningarTabOrder 
DesignSize�I  TLabelDDFakeFileEnabledLabelLeftTop-Width�Height;AnchorsakLeftakTopakRight AutoSizeCaption�   Tillåt direkta nedladdningar till vanliga lokala mappar (t.ex. Window Explorer). Tillåt inte nedladdningar till andra destinationer (ZIP-arkiv, FTP, etc.). Använd Dra && släpp skaltillägg, när det är tillgängligt.FocusControlDDFakeFileEnabledButtonWordWrap	OnClickDDLabelClick  TLabelDDFakeFileDisabledLabelLeftTop� Width�Height<AnchorsakLeftakTopakRight AutoSizeCaption�   Möjliggör nerladdningar till valfri destination (vanliga kataloger, ZIP-arkiv, FTP, etc.). Filer laddas först ner till en temporär katalog och flyttas därefter till destinationen.FocusControlDDFakeFileDisabledButtonWordWrap	OnClickDDLabelClick  TLabelDragExtStatusLabelLeftToplWidthdHeightCaptionDragExtStatusLabelFocusControlDDFakeFileEnabledButtonShowAccelCharOnClickDDLabelClick  TLabelDDDrivesLabelLeftTop~Width� HeightCaption7   Tillåt att filer släpps till dessa &nätverksenheter:FocusControlDDDrivesMemo  TRadioButtonDDFakeFileEnabledButtonLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption4   Bestäm mål för släpp genom att dra en &falsk filTabOrder OnClickControlChange  TRadioButtonDDFakeFileDisabledButtonLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption$   Ladda ner filer via tillfällig mappTabOrderOnClickControlChange  	TCheckBoxDDWarnLackOfTempSpaceCheckLeftTop.Width;HeightAnchorsakLeftakTopakRight Caption)   &Varna vid otillräckligt med diskutrymmeTabOrderOnClickControlChange  TMemoDDDrivesMemoLeftTop� Width�HeightBAnchorsakLeftakTopakRight Lines.StringsDDDrivesMemo 
ScrollBars
ssVerticalTabOrder    	TTabSheet
QueueSheetTagHelpType	htKeywordHelpKeywordui_pref_backgroundCaptionBakgrund
ImageIndex
TabVisible
DesignSize��  	TGroupBox
QueueGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Överföringar i bakgrundenTabOrder 
DesignSize��   TLabelLabel5Left	TopWidth� HeightCaption)   &Maximalt antal samtidiga överföringar:FocusControlQueueTransferLimitEdit  TLabelQueueKeepDoneItemsCheckLeftTop� Width� HeightCaption*   Visa avslutade överföringar i kön för:FocusControlQueueKeepDoneItemsForComboOnClickControlChange  TLabel"ParallelTransferThresholdUnitLabelLeft� Top� WidthHeightCaptionbyteFocusControlParallelTransferThresholdComboOnClickControlChange  TUpDownEditQueueTransferLimitEditLefteTopWidthOHeight	AlignmenttaRightJustifyMaxValue       �@MinValue       ��?AnchorsakTopakRight 	MaxLengthTabOrder   	TCheckBoxQueueAutoPopupCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight CaptionC   Visa bakgrundsöverföringarnas prompt &automatiskt vid inaktivitetTabOrder  	TCheckBox
QueueCheckLeftTopEWidth�HeightAnchorsakLeftakTopakRight Caption$   &Överför som standard i bakgrundenTabOrder  	TCheckBoxQueueNoConfirmationCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption1   I&ngen bekräftelser för bakgrundsöverföringarTabOrder  	TCheckBoxQueueParallelCheckLeftTop\Width�HeightAnchorsakLeftakTopakRight Caption3   &Använd flera anslutningar för enkel överföringTabOrderOnClickControlChange  	TCheckBoxEnableQueueByDefaultCheckLeftTop.Width�HeightAnchorsakLeftakTopakRight Caption$   &Aktivera köbehandling som standardTabOrder  	TComboBoxQueueKeepDoneItemsForComboLeftITop� WidthkHeightStylecsDropDownListAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeItems.StringsAldrig15 sekunder1 minut
15 minuter1 timmeAlltid   	TCheckBoxParallelTransferCheckLeftTopsWidth�HeightAnchorsakLeftakTopakRight Caption4   &Använd flera anslutningar för enstaka filer ovan:TabOrderOnClickControlChange  	TComboBoxParallelTransferThresholdComboLeft+Top� WidthfHeightAnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChangeOnExitSizeComboExitItems.Strings1M10M100M1G    	TGroupBoxQueueViewGroupLeftTop� Width�Height_AnchorsakLeftakTopakRight Caption   KölistaTabOrder
DesignSize�_  TRadioButtonQueueViewShowButtonLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionVi&saTabOrder   TRadioButtonQueueViewHideWhenEmptyButtonLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption   &Dölj ifall tomTabOrder  TRadioButtonQueueViewHideButtonLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption   &DöljTabOrder    	TTabSheetStorageSheetTagHelpType	htKeywordHelpKeywordui_pref_storageCaptionLagring
ImageIndex
TabVisible
DesignSize��  	TGroupBoxStorageGroupLeftTopWidth�Height`AnchorsakLeftakTopakRight Caption   Inställningar för lagringTabOrder 
DesignSize�`  
TPathLabelAutomaticIniFileStorageLabelLeft� Top-Width� HeightActiveTextColorclWindowTextIndentHorizontal IndentVertical InactiveTextColor
clGrayTextOnGetStatus%AutomaticIniFileStorageLabelGetStatusAlignalNoneAnchorsakLeftakTopakRight AutoSize  TRadioButtonRegistryStorageButtonLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionWindowsre&gistretTabOrder OnClickControlChange  TRadioButtonAutomaticIniFileStorageButtonLeftTop-Width� HeightCaption&Automatisk INI-filTabOrderOnClickControlChange  TRadioButtonCustomIniFileStorageButtonLeftTopDWidth� HeightCaptionA&npassad INI-filTabOrderOnClickCustomIniFileStorageButtonClick  TFilenameEditCustomIniFileStorageEditLeft� TopAWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialog#CustomIniFileStorageEditAfterDialog
DialogKinddkSave
DefaultExtiniFilter*INI-fil (*.ini)|*.ini|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist ClickKey@AnchorsakLeftakTopakRight TabOrderTextCustomIniFileStorageEditOnChangeControlChangeOnExitCustomIniFileStorageEditExit   	TGroupBoxTemporaryDirectoryGrouoLeftTophWidth�Height� AnchorsakLeftakTopakRight Caption   Temporär katalogTabOrder
DesignSize��   TLabelLabel6Left	TopWidth�HeightAnchorsakLeftakTopakRight AutoSizeCaption?   Ange var nerladdade och redigerade filer ska sparas temporärt.FocusControl DDSystemTemporaryDirectoryButtonShowAccelCharWordWrap	  TRadioButton DDSystemTemporaryDirectoryButtonLeftTop5Width�HeightAnchorsakLeftakTopakRight Caption%   &Använd systemets temporära katalogTabOrder OnClickControlChange  TRadioButton DDCustomTemporaryDirectoryButtonLeftTopLWidth� HeightCaption   Använd den här &katalogen:TabOrderOnClickControlChange  TDirectoryEditDDTemporaryDirectoryEditLeft� TopIWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogText2   Välj katalog för temporära dra && släpp filer.ClickKey@AnchorsakLeftakTopakRight TabOrderTextDDTemporaryDirectoryEditOnChangeControlChange  	TCheckBoxTemporaryDirectoryCleanupCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption.   &Rensa gamla temporära kataloger vid uppstartTabOrderOnClickControlChange  	TCheckBox%ConfirmTemporaryDirectoryCleanupCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption   &Fråga innan rensningTabOrderOnClickControlChange  	TCheckBox$TemporaryDirectoryAppendSessionCheckLeftTopcWidth�HeightAnchorsakLeftakTopakRight Caption3   Lägg till &sessionsnamn till temporära sökvägenTabOrderOnClickControlChange  	TCheckBox!TemporaryDirectoryAppendPathCheckLeftTopzWidth�HeightAnchorsakLeftakTopakRight Caption5   Lägg till f&järrsökväg till temporära sökvägenTabOrderOnClickControlChange  	TCheckBox$TemporaryDirectoryDeterministicCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight CaptionH   Behåll tillfälliga kopior av fjärrfiler i &deterministiska sökvägarTabOrderOnClickControlChange   	TGroupBoxOtherStorageGroupLeftTopFWidth�Height2AnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize�2  TLabelRandomSeedFileLabelLeft	TopWidth^HeightCaption   Sl&umptalsfröfil:FocusControlRandomSeedFileEdit  TFilenameEditRandomSeedFileEditLeft� TopWidth� HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPathEditAfterDialog
DialogKinddkSave
DefaultExtrndFilter4   Slumptalsfröfiler (*.rnd|*.rnd|Alla filer (*.*)|*.*DialogOptionsofHideReadOnlyofPathMustExist DialogTitle   Välj fil för slumptalsfröClickKey@AnchorsakLeftakTopakRight TabOrder TextRandomSeedFileEditOnChangeControlChange    	TTabSheetTransferEnduranceSheetTagHelpType	htKeywordHelpKeywordui_pref_resumeCaptionTolerans
ImageIndex
TabVisible
DesignSize��  	TGroupBox	ResumeBoxLeftTopWidth�Height|AnchorsakLeftakTopakRight Caption@   Aktivera överföringspaus/överför till temporär filnamn förTabOrder  TLabelResumeThresholdUnitLabel2Left}TopGWidthHeightCaptionKBFocusControlResumeThresholdEdit  TRadioButtonResumeOnButtonLeftTopWidth� HeightCaptionA&lla filerTabOrder OnClickControlChange  TRadioButtonResumeSmartButtonLeftTop-Width� HeightCaption   Filer stö&rre än:TabOrderOnClickControlChange  TRadioButtonResumeOffButtonLeftTopaWidth� HeightCaptionA&vaktiveraTabOrderOnClickControlChange  TUpDownEditResumeThresholdEditLeftTopDWidth\Height	AlignmenttaRightJustify	Increment       �@MaxValue       �@TabOrderOnClickControlChange   	TGroupBoxSessionReopenGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption   Automatisk återanslutningTabOrder
DesignSize��   TLabelSessionReopenAutoLabelLeftTop0WidthVHeightCaption   &Återanslut efter:FocusControlSessionReopenAutoEdit  TLabelSessionReopenAutoSecLabelLeftTop0Width+HeightCaptionsekunderFocusControlSessionReopenAutoEdit  TLabelSessionReopenTimeoutLabelLeft	Top� WidthxHeightCaption   &Fortsätt återansluta i:FocusControlSessionReopenTimeoutEdit  TLabelSessionReopenTimeoutSecLabelLeftTop� Width+HeightCaptionsekunderFocusControlSessionReopenTimeoutEdit  TLabelSessionReopenAutoStallLabelLeftTop� WidthVHeightCaption   Å&teranslut efter:FocusControlSessionReopenAutoStallEdit  TLabelSessionReopenAutoStallSecLabelLeftTop� Width+HeightCaptionsekunderFocusControlSessionReopenAutoStallEdit  TLabelSessionReopenAutoIdleLabelLeftTopdWidthVHeightCaption   Å&teranslut efter:FocusControlSessionReopenAutoIdleEdit  TLabelSessionReopenAutoIdleSecLabelLeftTopdWidth+HeightCaptionsekunderFocusControlSessionReopenAutoIdleEdit  	TCheckBoxSessionReopenAutoCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionA   &Automatiskt återanslut session, om den bryts under överföringTabOrder OnClickControlChange  TUpDownEditSessionReopenAutoEditLeft� Top-WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder  	TCheckBoxSessionReopenAutoIdleCheckLeftTopJWidth�HeightAnchorsakLeftakTopakRight Caption<   Automatiskt återanslut session, om den &bryts medan inaktivTabOrderOnClickControlChange  TUpDownEditSessionReopenTimeoutEditLeft� Top� WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue      ��@	MaxLengthTabOrder
OnGetValue SessionReopenTimeoutEditGetValue
OnSetValue SessionReopenTimeoutEditSetValue  	TCheckBoxSessionReopenAutoStallCheckLeftTop~Width�HeightAnchorsakLeftakTopakRight Caption0   Automatiskt återanslut session, om den &stannarTabOrderOnClickControlChange  TUpDownEditSessionReopenAutoStallEditLeft� Top� WidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder  TUpDownEditSessionReopenAutoIdleEditLeft� TopaWidthaHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��?Value       �@	MaxLengthTabOrder    	TTabSheetUpdatesSheetTagHelpType	htKeywordHelpKeywordui_pref_updatesCaptionUppdateringar
ImageIndex
TabVisible
DesignSize��  	TGroupBoxUpdatesGroup2LeftTopWidth�Height{AnchorsakLeftakTopakRight CaptionAutomatiska uppdateringarTabOrder 
DesignSize�{  TLabelLabel12Left	TopHWidth� HeightCaptionAutomatisk kontroll&period:FocusControlUpdatesPeriodCombo  TLabelUpdatesAuthenticationEmailLabelLeft	TopWidth� HeightCaption6   &E-postadress behörig för automatiska uppdateringar:FocusControlUpdatesAuthenticationEmailEdit  	TComboBoxUpdatesPeriodComboLeftFTopEWidthnHeightStylecsDropDownListAnchorsakTopakRight TabOrderItems.StringsAldrigDagligVeckovis
   Månadsvis   	TCheckBoxUpdatesShowOnStartupLeftTopbWidth�HeightAnchorsakLeftakTopakRight Caption-&Visa information om uppdatering vid uppstartTabOrderOnClickControlChange  TEditUpdatesAuthenticationEmailEditLeft	Top(Width8HeightAnchorsakLeftakTopakRight TabOrder OnChangeControlChangeOnExit"UpdatesAuthenticationEmailEditExit  TStaticTextUpdatesLinkLeftFTop,Width@HeightAnchorsakTopakRight Caption   Läs merTabOrderTabStop	OnClickUpdatesLinkClick   	TGroupBoxUpdatesProxyGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption
AnslutningTabOrder
DesignSize��   TLabelUpdatesProxyHostLabelLeftTop[Width[HeightCaption   Proxy &värdnamn:FocusControlUpdatesProxyHostEdit  TLabelUpdatesProxyPortLabelLeftFTop[WidthFHeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlUpdatesProxyPortEdit  TUpDownEditUpdatesProxyPortEditLeftFTopmWidthnHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrder  TEditUpdatesProxyHostEditLeftTopmWidth&HeightAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextUpdatesProxyHostEdit  TRadioButtonUpdatesProxyCheckLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption   A&nvänd proxyserverTabOrderOnClickControlChange  TRadioButtonUpdatesDirectCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionIngen &proxyTabOrder OnClickControlChange  TRadioButtonUpdatesAutoCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption)   Detektera &automatisk proxyinställningarTabOrderOnClickControlChange   	TGroupBoxUpdatesOptionsGroupLeftTop� Width�HeightRAnchorsakLeftakTopakRight Caption
AlternativTabOrder
DesignSize�R  TLabelUpdatesBetaVersionsLabelLeftTopWidth~HeightCaption+Kontrollera ifall det finns &betaversioner:FocusControlUpdatesBetaVersionsCombo  	TComboBoxUpdatesBetaVersionsComboLeftFTopWidthnHeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TCheckBoxCollectUsageCheckLeftTop4Width>HeightAnchorsakLeftakTopakRight Caption"   Tillåt &anonym användarstatistikTabOrderOnClickControlChange  TButtonUsageViewButtonLeftFTop0WidthnHeightAnchorsakTopakRight CaptionVisa &statistikTabOrderOnClickUsageViewButtonClick    	TTabSheetCopyParamListSheetTagHelpType	htKeywordHelpKeywordui_pref_transferCaption	   Överför
ImageIndex
TabVisible
DesignSize��  	TGroupBoxCopyParamListGroupLeftTopWidth�Height�AnchorsakLeftakTopakRightakBottom Caption   Överför förinställningarTabOrder 
DesignSize��  TLabelCopyParamLabelLeft	TopFWidth�Height5AnchorsakLeftakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamLabelClick  	TListViewCopyParamListViewLeft	TopWidth�Height*AnchorsakLeftakTopakRightakBottom ColumnsCaption   Beskrivning förinställningarWidthd Caption
AutomatiskWidth(  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder 	ViewStylevsReportOnCustomDrawItemCopyParamListViewCustomDrawItemOnDataCopyParamListViewData
OnDblClickCopyParamListViewDblClick	OnEndDragListViewEndDrag
OnDragDropCopyParamListViewDragDrop
OnDragOverCopyParamListViewDragOver	OnKeyDownCopyParamListViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddCopyParamButtonLeft	Top~WidthZHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddCopyParamButtonClick  TButtonRemoveCopyParamButtonLeft	Top�WidthZHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveCopyParamButtonClick  TButtonUpCopyParamButtonLeftZTop~WidthZHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownCopyParamButtonClick  TButtonDownCopyParamButtonLeftZTop�WidthZHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownCopyParamButtonClick  TButtonEditCopyParamButtonLeftiTop~WidthZHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickEditCopyParamButtonClick  TButtonDuplicateCopyParamButtonLeftiTop�WidthZHeightAnchorsakLeftakBottom Caption&Dubblera...TabOrderOnClickDuplicateCopyParamButtonClick  	TCheckBoxCopyParamAutoSelectNoticeCheckLeftTop�Width�HeightAnchorsakLeftakRightakBottom CaptionS   &Meddela när överföringsinställningarna automatiskt använder de förinställdaTabOrderOnClickControlChange    	TTabSheetWindowSheetTagHelpType	htKeywordHelpKeywordui_pref_windowCaption   Fönster
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPathInCaptionGroupLeftTopWidth�Height_AnchorsakLeftakTopakRight Caption   Sökväg i fönstertitelTabOrder
DesignSize�_  TRadioButtonPathInCaptionFullButtonLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Visa &lång sökvägTabOrder   TRadioButtonPathInCaptionShortButtonLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption   Visa &kort sökvägTabOrder  TRadioButtonPathInCaptionNoneButtonLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption
Visa &inteTabOrder   	TGroupBoxWindowMiscellaneousGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption   ÖvrigtTabOrder
DesignSize��   	TCheckBoxMinimizeToTrayCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionN   &Minimera huvudfönstret till aktivitetsfältets statusområde (systemfältet)TabOrder OnClickControlChange  	TCheckBox&ExternalSessionInExistingInstanceCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption>   Öppna nya externa initierade sessioner i &befintliga fönsterTabOrderOnClickControlChange  	TCheckBoxKeepOpenWhenNoSessionCheckLeftTop[Width�HeightAnchorsakLeftakTopakRight CaptionA   &Håll huvudfönstret öppet när den sista sessionen är stängdTabOrderOnClickControlChange  	TCheckBoxShowTipsCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption&Visa tips vid uppstartTabOrderOnClickControlChange  	TCheckBoxShowLoginWhenNoSessionCheckLeftTopDWidth�HeightAnchorsakLeftakTopakRight CaptionO   &Visa inloggningsdialogrutan vid start och när den sista sessionen är stängdTabOrderOnClickControlChange  	TCheckBox SessionTabCaptionTruncationCheckLeftToprWidth�HeightAnchorsakLeftakTopakRight Caption4   &Trunkera fliktitlar när de inte passar i fönstretTabOrderOnClickControlChange   	TGroupBoxWorkspacesGroupLeftTopWidth�HeightwAnchorsakLeftakTopakRight Caption
ArbetsytorTabOrder 
DesignSize�w  TLabelAutoWorkspaceLabelLeftTop-Width� HeightCaption&Standardnamn arbetsyta:FocusControlAutoWorkspaceCombo  	TCheckBoxAutoSaveWorkspaceCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption'Spara &automatiskt arbetsyta vid avslutTabOrder OnClickControlChange  	TComboBoxAutoWorkspaceComboLeftTop?Width�HeightAnchorsakLeftakTopakRight DropDownCountTabOrderOnClickControlChange  	TCheckBoxAutoSaveWorkspacePasswordsCheckLeftTop\Width�HeightAnchorsakLeftakTopakRight Caption#Save &passwords (not recommended) XTabOrderOnClickControlChange    	TTabSheetSecuritySheetTagHelpType	htKeywordHelpKeywordui_pref_securityCaption	   Säkerhet
ImageIndex
TabVisible
DesignSize��  	TGroupBoxMasterPasswordGroupLeftTopWidth�HeightPAnchorsakLeftakTopakRight Caption   HuvudlösenordTabOrder 
DesignSize�P  TButtonSetMasterPasswordButtonLeft	Top-WidthHeightCaption   Ä&ndra huvudlösenord...TabOrderOnClickSetMasterPasswordButtonClick  	TCheckBoxUseMasterPasswordCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   An&vänd huvudlösenordTabOrder OnClickUseMasterPasswordCheckClick   	TGroupBoxPasswordGroupBoxLeftTopXWidth�Height0AnchorsakLeftakTopakRight Caption   SessionslösenordTabOrder
DesignSize�0  	TCheckBoxSessionRememberPasswordCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption1   Kom ihåg &lösenord under sessionens varaktighetTabOrder    	TGroupBoxSshHostCAsGroupLeftTop� Width�HeightKAnchorsakLeftakTopakRightakBottom Caption"   Betrodda värdcertifikatutfärdareTabOrder
DesignSize�K  	TListViewSshHostCAsViewLeft	Top-Width�Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionNamnWidthd Caption   VärdarWidthd  ColumnClickDoubleBuffered	HideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedTabOrder	ViewStylevsReportOnDataSshHostCAsViewData
OnDblClickSshHostCAsViewDblClick	OnKeyDownSshHostCAsViewKeyDownOnSelectItemListViewSelectItem  TButtonAddSshHostCAButtonLeft	Top(WidthZHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddSshHostCAButtonClick  TButtonRemoveSshHostCAButtonLeft� Top(WidthZHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveSshHostCAButtonClick  TButtonEditSshHostCAButtonLeftiTop(WidthZHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickEditSshHostCAButtonClick  	TCheckBoxSshHostCAsFromPuTTYCheckLeftTopWidth�HeightCaption    &Ladda behörigheter från PuTTYTabOrder OnClickSshHostCAsFromPuTTYCheckClick  TButtonConfigureSshHostCAsButtonLeft	Top(Width� HeightAnchorsakLeftakBottom Caption&Redigera i PuTTY...TabOrderOnClickConfigureSshHostCAsButtonClick    	TTabSheetIntegrationAppSheetTagHelpType	htKeywordHelpKeywordui_pref_integration_appCaptionApplikationer
ImageIndex
TabVisible
DesignSize��  	TGroupBoxExternalAppsGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionExterna applikationerTabOrder 
DesignSize��   TLabelPuttyPathLabelLeft	TopWidth� HeightCaption    &PuTTY/Terminal klient sökväg:FocusControlPuttyPathEdit  TLabelPuttyRegistryStorageKeyLabelLeft	Top� WidtheHeightCaptionPuTTY registernyc&kelFocusControlPuttyRegistryStorageKeyEdit  THistoryComboBoxPuttyPathEditLeft	Top(WidthUHeightAnchorsakLeftakTopakRight TabOrder OnChangePuttyPathEditChangeOnExitPuttyPathEditExit  	TCheckBoxPuttyPasswordCheck2LeftTopUWidth�HeightAnchorsakLeftakTopakRight Caption?   &Kom ihåg sessionslösenord och överför det till PuTTY (SSH)TabOrder  	TCheckBoxAutoOpenInPuttyCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption)   &Öppna automatiskt en ny session i PuTTYTabOrder  TButtonPuttyPathBrowseButtonLeftdTop'WidthPHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClickPuttyPathBrowseButtonClick  	TCheckBoxTelnetForFtpInPuttyCheckLeftToplWidth�HeightAnchorsakLeftakTopakRight Caption2   Öppna &Telnetsessioner i PuTTY för FTP-sessionerTabOrder  TStaticTextPuttyPathHintTextLeft� Top?Width~Height	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	   &mönsterTabOrderTabStop	  THistoryComboBoxPuttyRegistryStorageKeyEditLeft	Top� Width�HeightStylecsDropDownListAnchorsakLeftakTopakRight TabOrderOnChangeControlChange    	TTabSheetNetworkSheetTagHelpType	htKeywordHelpKeywordui_pref_networkCaption   Nätverk
ImageIndex
TabVisible
DesignSize��  	TGroupBoxExternalIpAddressGroupBox2LeftTopWidth�Height� AnchorsakLeftakTopakRight Caption*   Inkommande FTP-anslutningar (aktivt läge)TabOrder 
DesignSize��   TLabelLocalPortNumberRangeLabelLeft|TopzWidthHeightCaption      TRadioButtonRetrieveExternalIpAddressButtonLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption/   Hämta extern IP-adress från &operativsystemetTabOrder OnClickControlChange  TRadioButtonCustomExternalIpAddressButtonLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption%   Använd &följande externa IP-adress:TabOrderOnClickControlChange  TEditCustomExternalIpAddressEditLeftTopCWidth� HeightTabOrderOnClickControlChange  	TCheckBoxLocalPortNumberCheckLeftTop`Width�HeightAnchorsakLeftakTopakRight Caption    Begränsa lyssnings&portar till:TabOrderOnClickControlChange  TUpDownEditLocalPortNumberMinEditLeftTopwWidth[Height	AlignmenttaRightJustifyMaxValue      ��@MinValue       �	@TabOrderOnChangeControlChangeOnExitLocalPortNumberMinEditExit  TUpDownEditLocalPortNumberMaxEditLeft� TopwWidth[Height	AlignmenttaRightJustifyMaxValue      ��@MinValue       �	@TabOrderOnChangeControlChangeOnExitLocalPortNumberMaxEditExit   	TGroupBoxConnectionsGroupLeftTop� Width�Height1AnchorsakLeftakTopakRight CaptionAnslutningarTabOrder
DesignSize�1  	TCheckBoxTryFtpWhenSshFailsCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption-   När SFTP-anslutning av&visas, portknacka FTPTabOrder OnClickControlChange    	TTabSheetPanelRemoteSheetTagHelpType	htKeywordHelpKeywordui_pref_panels_remoteCaption   Fjärr
ImageIndex
TabVisible
DesignSize��  	TGroupBoxPanelsRemoteDirectoryGroupLeftTopWidth�HeightbAnchorsakLeftakTopakRight Caption   FjärrpanelTabOrder 
DesignSize�b  TLabelRefreshRemoteDirectoryUnitLabelLeft�TopDWidthHeightAnchorsakTopakRight CaptionsShowAccelChar  	TCheckBoxShowInaccesibleDirectoriesCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Vis&a oåtkomliga katalogerTabOrder OnClickControlChange  	TCheckBoxAutoReadDirectoryAfterOpCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption:Uppdatera auto&matisk katalog efter operation (CTRL+ALT+R)TabOrderOnClickControlChange  	TCheckBoxRefreshRemotePanelCheckLeftTopDWidthBHeightAnchorsakLeftakTopakRight Caption   Uppdatera fjärrpanel varj&eTabOrderOnClickControlChange  TUpDownEditRefreshRemotePanelIntervalEditLeftWTopAWidthQHeight	AlignmenttaRightJustify	Increment       �@MaxValue      <�@MinValue       �@AnchorsakTopakRight 	MaxLengthTabOrderOnChangeControlChange    	TTabSheetPanelLocalSheetTagHelpType	htKeywordHelpKeywordui_pref_panels_localCaptionLokal
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLocalPanelGroupLeftTopWidth�Height_AnchorsakLeftakTopakRight CaptionLokal panelTabOrder 
DesignSize�_  	TCheckBoxPreserveLocalDirectoryCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption/   &Ändra inte tillstånd när du byter sessionerTabOrderOnClickControlChange  	TCheckBoxSystemContextMenuCheckLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption   Använd filsystemets snabbmenyTabOrderOnClickControlChange  	TCheckBoxDeleteToRecycleBinCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption!&Ta bort filer till papperskorgenTabOrder OnClickControlChange    	TTabSheetLanguagesSheetTagCaption   Språk
ImageIndex
TabVisible
DesignSize��  	TGroupBoxLanguagesGroupLeftTopWidth�Height�AnchorsakLeftakTopakRightakBottom Caption   SpråkTabOrder 
DesignSize��  TLabelLanguageChangeLabelLeft	Top�Width� HeightAnchorsakLeftakBottom Caption-   Ändringar börjar gälla efter nästa start.ShowAccelChar  	TListViewLanguagesViewLeft	TopWidth�Height�AnchorsakLeftakTopakRightakBottom ColumnsAutoSize	  DoubleBuffered	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedShowColumnHeadersTabOrder 	ViewStylevsReportOnCustomDrawItemLanguagesViewCustomDrawItemOnSelectItemListViewSelectItem  TButtonLanguagesGetMoreButtonLeftFTop�WidthnHeightAnchorsakRightakBottom Caption   Hämta &fler...TabOrderOnClickLanguagesGetMoreButtonClick    	TTabSheetEditorInternalSheetTagHelpType	htKeywordHelpKeywordui_pref_editor_internalCaptionIntern editor
TabVisible
DesignSize��  	TGroupBoxInternalEditorGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionVisningTabOrder 
DesignSize��   TLabelLabel9Left	Top-WidthKHeightCaption&Tabulatorstorlek:FocusControlEditorTabSizeEdit  TLabelLabel11Left	Top\Width^HeightCaptionStandard&kodning:FocusControlEditorEncodingCombo  	TCheckBoxEditorWordWrapCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Ko&rta av långa raderTabOrder OnClickControlChange  TUpDownEditEditorTabSizeEditLeft	Top?Width� Height	AlignmenttaRightJustifyMaxValue       �@MinValue       ��?	MaxLengthTabOrderOnChangeControlChange  	TComboBoxEditorEncodingComboLeft	TopnWidth� HeightStylecsDropDownList	MaxLengthTabOrderOnChangeControlChange   	TGroupBox	FontGroupLeftTop� Width�HeightwAnchorsakLeftakTopakRight CaptionFontTabOrder
DesignSize�w  TLabelEditorFontLabelLeft� TopWidthHeightWAnchorsakLeftakTopakRightakBottom AutoSizeCaptionEditorFontLabelColorclWhiteParentColorShowAccelCharTransparent
OnDblClickEditorFontLabelDblClick  TButtonEditorFontButtonLeft	TopWidth� HeightCaption   &Välj font...TabOrder OnClickEditorFontButtonClick  TButtonEditorFontColorButtonLeft	Top5Width� HeightCaption
   &TextfärgTabOrderOnClickEditorFontColorButtonClick  TButtonEditorBackgroundColorButtonLeft	TopTWidth� HeightCaptionStandard&bakgrundTabOrderOnClick EditorBackgroundColorButtonClick   	TGroupBoxInternalEditorBehaviourGroupLeftTopWidth�Height1AnchorsakLeftakTopakRight CaptionBeteendeTabOrder
DesignSize�1  	TCheckBoxEditorDisableSmoothScrollCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Inaktivera &jämn rullningTabOrder OnClickControlChange    	TTabSheetFileColorsSheetTagHelpType	htKeywordHelpKeywordui_pref_file_colorsCaption
   Filfärger
ImageIndex
TabVisible
DesignSize��  	TGroupBoxFileColorsGroupLeftTopWidth�Height�AnchorsakLeftakTopakRightakBottom Caption
   FilfärgerTabOrder 
DesignSize��  	TListViewFileColorsViewLeft	TopWidth�HeightyAnchorsakLeftakTopakRightakBottom Columns  ColumnClickDoubleBuffered	DragModedmAutomaticHideSelection	OwnerData	ReadOnly		RowSelect	ParentDoubleBufferedParentShowHintShowColumnHeadersShowHintTabOrder 	ViewStylevsReportOnCustomDrawItemFileColorsViewCustomDrawItemOnDataFileColorsViewData
OnDblClickFileColorsViewDblClick	OnEndDragListViewEndDrag
OnDragDropFileColorsViewDragDrop
OnDragOverListViewDragOver	OnKeyDownFileColorsViewKeyDownOnSelectItemListViewSelectItemOnStartDragListViewStartDrag  TButtonAddFileColorButtonLeft	Top�WidthZHeightAnchorsakLeftakBottom Caption   &Lägg till...TabOrderOnClickAddEditFileColorButtonClick  TButtonRemoveFileColorButtonLeft	Top�WidthZHeightAnchorsakLeftakBottom Caption&Ta bortTabOrderOnClickRemoveFileColorButtonClick  TButtonUpFileColorButtonLeftZTop�WidthZHeightAnchorsakRightakBottom Caption&UppTabOrderOnClickUpDownFileColorButtonClick  TButtonDownFileColorButtonLeftZTop�WidthZHeightAnchorsakRightakBottom Caption&NerTabOrderOnClickUpDownFileColorButtonClick  TButtonEditFileColorButtonLeftiTop�WidthZHeightAnchorsakLeftakBottom Caption&Redigera...TabOrderOnClickAddEditFileColorButtonClick    	TTabSheetSearchSheetHelpType	htKeywordHelpKeywordui_pref_searchCaptionSearchSheet
ImageIndex
TabVisible
DesignSize��  	TGroupBoxSearchGroupLeftTopWidth�Height�AnchorsakLeftakTopakRightakBottom Caption   SökTabOrder     TPanel	LeftPanelLeft Top Width� Height�AlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� �  TPanelNavigationPanelLeftTop$Width� Height�AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder 	TTreeViewNavigationTreeLeft Top Width� Height�AlignalClientDoubleBuffered	HideSelectionHotTrack	IndentParentDoubleBufferedReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChange
OnChangingNavigationTreeChangingOnCollapsingNavigationTreeCollapsingOnEnterNavigationTreeEnterItems.NodeData
�     6          ��������           E n v i r o n m e n t X 2          ��������            
I n t e r f a c e X ,          ��������            W i n d o w X 2          ��������            
C o m m a n d e r X 0          ��������            	E x p l o r e r X 2          ��������            
L a n g u a g e s X ,          ��������           P a n e l s X 6          ��������            F i l e   c o l o r s X ,          ��������            R e m o t e X *          ��������            L o c a l X ,          ��������           E d i t o r X >          ��������            I n t e r n a l   e d i t o r X 0          ��������           	T r a n s f e r X 0          ��������            	D r a g D r o p X 4          ��������            B a c k g r o u n d X ,          ��������            R e s u m e X .          ��������            N e t w o r k X 0          ��������            	S e c u r i t y X .          ��������            L o g g i n g X 6       	   ��������           I n t e g r a t i o n X 8          ��������            A p p l i c a t i o n s X 0       
   ��������            	C o m m a n d s X .          ��������            S t o r a g e X .          ��������            U p d a t e s X    
TComboEdit
SearchEditLeftTopWidth� HeightHelpType	htKeywordHelpKeywordui_pref_searchButtonTabStopButtonCaption   'ClickKey AnchorsakLeftakTopakRight TabOrder OnButtonClickSearchEditButtonClickOnChangeSearchEditChangeEnterOnEnterSearchEditChangeEnter    TButton
HelpButtonLeftTop�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelComponentsPanelLeft TopWidth]Height2AlignalBottom
BevelOuterbvNoneColorclWindowParentBackgroundTabOrder  
TPopupMenuRegisterAsUrlHandlerMenuLeft8Top� 	TMenuItemRegisterAsUrlHandlerItemCaption
RegistreraOnClickRegisterAsUrlHandlerItemClick  	TMenuItemMakeDefaultHandlerItemCaption   Gör WinSCP &standardprogram...OnClickMakeDefaultHandlerItemClick  	TMenuItem!UnregisterForDefaultProtocolsItemCaptionAvregistreraOnClick&UnregisterForDefaultProtocolsItemClick   
TPopupMenuAddCommandMenuLeft� Top� 	TMenuItemAddCustomCommandMenuItemCaption    Lägg till &anpassat kommando...OnClickAddCustomCommandMenuItemClick  	TMenuItemAddExtensionMenuItemCaption   Lägg till &utökning...OnClickAddExtensionMenuItemClick      TPF0TProgressFormProgressFormLeft�Top#HelpType	htKeywordHelpKeywordui_progressBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption	OperationClientHeight&ClientWidth�ColorclWindowFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 	PopupModepmAutoPositionpoOwnerFormCenterOnHideFormHideOnShowFormShow
DesignSize�& 
TextHeight 	TPaintBoxAnimationPaintBoxLeftTopWidth Height   TPanel	MainPanelLeft2TopWidthTHeightEAnchorsakLeftakTopakRight 
BevelOuterbvNoneParentColor	TabOrder 
DesignSizeTE  TLabel	PathLabelLeft TopWidthHeightCaptionFileX:ShowAccelChar  
TPathLabel	FileLabelLeft8TopWidthHeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelTargetLabelLeft TopWidth$HeightCaption   Mål:ShowAccelChar  
TPathLabelTargetPathLabelLeft8TopWidthHeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TProgressBarOperationProgressLeft Top+WidthTHeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder    TPanelTransferPanelLeft2TopLWidthhHeight@AnchorsakLeftakTopakRight 
BevelOuterbvNoneParentColor	TabOrder
DesignSizeh@  TLabelStartTimeLabelLefthTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00ShowAccelChar  TLabelTimeLeftLabelLefthTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption00:00:00ShowAccelChar  TLabelTimeLeftLabelLabelLeft TopWidth2HeightCaption	Tid kvar:ShowAccelChar  TLabelCPSLabelLeft
TopWidthJHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption0 KB/sShowAccelChar  TLabelTimeElapsedLabelLeft
TopWidthJHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption00:00:00ShowAccelChar  TLabelBytesTransferredLabelLefthTopWidthAHeight	AlignmenttaRightJustifyAutoSizeCaption0 KBShowAccelChar  TLabelLabel3Left� TopWidthIHeightAnchorsakTopakRight Caption   Förfluten tid:ShowAccelChar  TLabelStartTimeLabelLabelLeft TopWidth6HeightCaption
Start tid:ShowAccelChar  TLabelLabel4Left TopWidth[HeightCaption   Bytes överförda:ShowAccelChar  TLabelLabel12Left� TopWidth#HeightAnchorsakTopakRight Caption
Hastighet:ShowAccelChar  TProgressBarFileProgressLeft Top&WidthTHeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder    TPanelToolbarPanelLeft2Top� Width.HeightAnchorsakLeftakBottom 
BevelOuterbvNoneParentColor	TabOrder TTBXDockDockLeft Top Width.Height	AllowDragColorclWindow TTBXToolbarToolbarLeft Top DockModedmCannotFloatOrChangeDocksDragHandleStyledhNoneImages	ImageListParentShowHintProcessShortCuts	ShowHint	TabOrder ColorclWindow TTBXItem
CancelItemCaption&CancelX
ImageIndex ShortCutOnClickCancelItemClick  TTBXItemSkipItemCaption   &Hoppa över den här filen
ImageIndex	OnClickSkipItemClick  TTBXItemMinimizeItemCaption	&Minimera
ImageIndexShortCutM�  OnClickMinimizeItemClick  TTBXItemMoveToQueueItemCaption   Fortsätt i &bakgrunden
ImageIndexShortCutB�  OnClickMoveToQueueItemClick  TTBXSubmenuItemCycleOnceDoneItemCaption   När operationen är klarDropdownCombo	Hint3   Åtgärd som ska utföras när operationen är klar
ImageIndexShortCutF�  OnClickCycleOnceDoneItemClick TTBXItemIdleOnceDoneItemCaption   &Förbli inaktivChecked	
ImageIndex	RadioItem	OnClickOnceDoneItemClick  TTBXItemDisconnectOnceDoneItemCaption   &Koppla ifrån session
ImageIndex	RadioItem	OnClickOnceDoneItemClick  TTBXItemSuspendOnceDoneItemCaption   &Försätt datorn i viloläge
ImageIndex	RadioItem	OnClickOnceDoneItemClick  TTBXItemShutDownOnceDoneItemCaption   &Stäng av datorn
ImageIndex	RadioItem	OnClickOnceDoneItemClick   TTBXComboBoxItemSpeedComboBoxItem	EditWidthnHint   Hastighetsbegränsning (kB/s)
ImageIndexShortCutS�  OnAcceptTextSpeedComboBoxItemAcceptTextOnClickSpeedComboBoxItemClick	ShowImage	OnAdjustImageIndex!SpeedComboBoxItemAdjustImageIndexOnItemClickSpeedComboBoxItemItemClick     TPanelComponentsPanelLeft Top� Width�HeightnAlignalBottom
BevelEdgesbeTop 	BevelKindbkFlat
BevelOuterbvNoneTabOrder  TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeft(Top�   TPngImageList	ImageList	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:34+01:00" xmp:MetadataDate="2022-09-01T10:57:34+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:180c2c88-0c60-ab4a-b417-9c9f76a6e069" xmpMM:DocumentID="adobe:docid:photoshop:b1118248-b8f9-3348-b679-1d9529e70ef5" xmpMM:OriginalDocumentID="xmp.did:d542fc81-8626-f34b-9a93-59aa7ca76804"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d542fc81-8626-f34b-9a93-59aa7ca76804" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:180c2c88-0c60-ab4a-b417-9c9f76a6e069" stEvt:when="2022-09-01T10:57:34+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�sa  ~IDATxڥ�=K�@��Kb� �"Zď�~D��ͥ]t�{��\�C���Gd��"�`t�"�����K��6ѡ!p���CDXf1-�o{N��H�Zի~���X���_Q�<�~�F�v��ӿJ�*ND�z��6��Y�vnBaË�}*�CT!�rA2��@�n�=0�ζ88��&�Dm,)�k��as�^Z��"	���I,����j
����F!HB���Iʖ����3���q�fN��(����:2@<xZ�Rލ�K��u� �n#��I�'�_�"8���d��8�י�ۑ�$�^c���m$���Kl3� ��C��kcӧ3�2x*q�%�@�ۿ��F��tͫ8nӨ5��ɱ˩�T��1{Lˬ��y�ήO�    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
B  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:49+01:00" xmp:MetadataDate="2022-09-01T11:07:49+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c268d7f3-d2fb-104b-a1d0-bb0a4d3ff770" xmpMM:DocumentID="adobe:docid:photoshop:2f11441a-416e-0c44-a239-1906973e411c" xmpMM:OriginalDocumentID="xmp.did:f4e92379-e79c-1e49-9b59-46651bc855c3"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:f4e92379-e79c-1e49-9b59-46651bc855c3" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c268d7f3-d2fb-104b-a1d0-bb0a4d3ff770" stEvt:when="2022-09-01T11:07:49+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����   IDATx�cd�0�0H�O��0�a0j �  O����.    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:21+01:00" xmp:MetadataDate="2022-09-01T11:07:21+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8d79b445-e579-aa4e-a511-7e6ea5d0f336" xmpMM:DocumentID="adobe:docid:photoshop:112a4d25-3396-0146-a130-67964781a8f7" xmpMM:OriginalDocumentID="xmp.did:42dd8fde-1e56-f54f-a1ad-43e2df677ddd"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:42dd8fde-1e56-f54f-a1ad-43e2df677ddd" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8d79b445-e579-aa4e-a511-7e6ea5d0f336" stEvt:when="2022-09-01T11:07:21+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>k�K  �IDATx�}�]HSa�����|:u�����-ݔ� *��袠���.���� �.r^楤t�X��M�tS�(h���n��:�9��9�VS��<�}y9�������Gx��5�:%��}D"�i�E&��nձE�����Nb�V֊n^��i��U�R.cdͨ��ǧ/��`��F�
! �8f��Z�;05��mbr"�oc%��?|�/���jI�(���������[H�Y�V����x><^Z-O�İ���u�8��;i��ձ���Mŀ�Cj��D��Olg[��C����h�*�[Ҳ���� e^Y��s�x�#cx}ćh&��S�؄aA�e}���qY�g�.t=x3��|��,/M,µ�e����$E��=��%�>���7�!�n���o�Qp��Γ_L/���j�Q"G�ܥ�	���?���0>O-���q�s:��H��z'�Jq�}4~
��A�[�֣B�R�j���g$�R��:&�&�9��M�`R�֪�R�1Rd�@��2\�I���d������{k�8`�8շ#�j�=���{kb��t��
����r�V�[��� ��|#{���!W*9��*���8��i�56�8�-`�Q�]�ݪ���e�Ǳ��� �jM-K�	�    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:25+01:00" xmp:MetadataDate="2022-09-01T11:07:25+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c81b4c70-3613-134b-a7e2-f7aeded61170" xmpMM:DocumentID="adobe:docid:photoshop:c6dc1ac0-908a-694a-816e-ebaf60abec42" xmpMM:OriginalDocumentID="xmp.did:dfd8d9a0-d1be-f34f-9d41-200adc72f0d4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:dfd8d9a0-d1be-f34f-9d41-200adc72f0d4" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c81b4c70-3613-134b-a7e2-f7aeded61170" stEvt:when="2022-09-01T11:07:25+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>N
�   �IDATxڅ�_HSQ���m��6�F��Vsw�V�
�K(��&A�FT�=�>������A
!��^�N%Et:�j������mw���a65�q~�p~�������ض�a���ׁ�H�"����"����$�>��ӑg�Z���I�t�EA��D��LJN+��(�]�q��^@�f��7M�q�h1UXt(�v���������3Aء�m����$�[\��a��?���zRJ+���j�� <os;��tH��c���	�|^�X2>7�x��x)�դX�qPvĪ�9��Y��tއ� � 2�����:b���J
�F/�c�`��vC(���/Ky�r�ݒ�����,�����^��"���#��
-���a�#��6�*���>U����q!%�>QC ��YG�=j��.S��ne����8|�ġ�����OԎ�ou���`|�Xƪc3Z���(v����h���A��N�c�^���'�Y��sG������j�i$�Zĩ�1
�bEdI�'��tij�i�jxk��42�8�'R�3BJZ���@1��(�eY���gv]n䰛a��|�[�&��?�|��f0P~�C�Fג+�D�	��]�SL��6�]�$9Q�^&I���
90Q�YȚ�z�K&�7�P�����8�+*L�7��?
B��*�;N���(�[��UՖ),    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:30+01:00" xmp:MetadataDate="2022-09-01T11:07:30+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0091a1ba-ca2b-2540-8058-0145f5097785" xmpMM:DocumentID="adobe:docid:photoshop:517d3f28-5032-4548-b484-e16684345bec" xmpMM:OriginalDocumentID="xmp.did:365a17c0-743d-0d40-bf23-62e182bd42a2"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:365a17c0-743d-0d40-bf23-62e182bd42a2" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0091a1ba-ca2b-2540-8058-0145f5097785" stEvt:when="2022-09-01T11:07:30+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>m�$�  �IDATx�}�iHTQ��o��7�m��}T+�4B""�A4hC-���"#3(?�J"���dˇ����(jcj3�㘚��7����H��9����s��VҠ��ΣH"O�LFEI|1j��DI����j�j�E� �[ɒ
�(�������&���97qb+@�9�ݧ֪���r
��;@Icl��%�q�8��"��7_�F������8w����;���3��T8z)�b �m�G��@)�bȧ!9��c��0�l�$��O��x��y��� �����AQ�/��,xo��( ���6rq7��gU��
i�,j�BCQh�
�
���1Y,A����6�7=C��1d�5x`��'ˢ���@O�x�����Dz�ghX��ll�U�����D�!��Z%{+B��zo����M(������?{�kc�`|v�ru5em�Q1�
w:L����H��{�܏Q�-Ǎ�x��݇���#����ڂj�t|�O/C��
"�VQ,ȵ��W���/���a5#�~�:�~a�{ڊ�t+�a�ã�H
� !�T}S�\�912PD�;+Lg���3�2�;XG�v�@��ג�^�@�ac'�@�Tݍ�C��m���1��z�%Q�e�Pť��m��������h���2�.�՝Υ��E�jL�S./�X\J��Bi��)5{�	���Ƈg���*��� ��Q���a�    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:28+01:00" xmp:MetadataDate="2022-09-01T11:07:28+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0b476a77-d74a-3a4c-ab52-304f230a90f8" xmpMM:DocumentID="adobe:docid:photoshop:4cfee566-e453-214c-8355-090c9aea2e55" xmpMM:OriginalDocumentID="xmp.did:8423c53f-c864-744c-86c2-0a711a30412a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8423c53f-c864-744c-86c2-0a711a30412a" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0b476a77-d74a-3a4c-ab52-304f230a90f8" stEvt:when="2022-09-01T11:07:28+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  cIDATx�cd���Ul
���L���1(�|9���	��g`p�NO>`�s�I�r2 biA6.&V&��+RcQtϙ��������?<a�0�lVRS��)Į�!�����N�z����w�¨��R67S�$'L3�i�!�4� 2
�d�'�2*-�t�W�S����D��<��t� `dTZz��7;��fθ}��(���'�Ů���`#��0��;ff����t���7�D9�B���������肧[ր�1{>�ɓ'n޸����~~��fV���tFp �p0vq
�q)�2��	�m�>kC\t8CbR
��r�,rb-�<|��=�0��'�=��	�FU���<,��L��*���ۖ,f8v�(É�� 	���ar����*��\�����{����|���Q������	#;�޾��[MQ�a��x0���>ɋ�0�$e%�&f�,���� !��0������peG>$M��Ǡ�:�#���q�VU�s�����{�?���-�6�ր� ))).N��@EVy������-C߼����=���g�����C80"T�	�60�����g�~  �����PB    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
@	  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:34+01:00" xmp:MetadataDate="2022-09-01T11:07:34+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8fa9e7d5-fe22-1c4f-a15e-a98105fdc327" xmpMM:DocumentID="adobe:docid:photoshop:6a1ab271-94bc-fb4c-b40b-b15058f12d21" xmpMM:OriginalDocumentID="xmp.did:cbc7d4bd-e57e-5f47-bad5-43889c99a346"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cbc7d4bd-e57e-5f47-bad5-43889c99a346" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8fa9e7d5-fe22-1c4f-a15e-a98105fdc327" stEvt:when="2022-09-01T11:07:34+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>)��6  IDATx�]�kHQ��3���qz�7�}�jJ�)��$���fT��"� �!&V�m�=�w�������>�k�*)��cwggv�Nw'�w�0s����?�0X��f昖G�+X��!���3�J1Ay1��7�::���g�_�f�RoLjd�8Ϛ��hX��bD1�X�sOH��;y���Ȑ�rppPX �ĉ放$�)�d�E#~�����dn��U��|�n���_��B`�/lJN��9���l� `�@"�>C��2P����"�r>�h{Z�dd�0hc���/��t٠F�V(��!E�!I��{�sԃ{{*����F��1;sw_/*�-�ֶ0���$��yV��FP=�H���Ձ�i�o֟ �]7�]�Ec���k�Gkhؑny���t��OH@A~R�-D��G�@x��P{�u������^>�R�C�!����|OU�`l|����|*�R�x�e!��E��w�?�}�J��e o��/�����V�N��ǎ,��9����]EŃ׼�B��Ck�N�hQ�$�aT�B�E�H������ <U-8��}\6Ѻ+��8��a�	�c���wQf���kj�n-z6W���M��Q1Q�ͶBM��Fp�bpqً����K����U-��oƗ&7���l*�:�U-,3�����~�����а�����d���&K_�ސRz�D��s<\Z<-ߝ�&��r-��<$�`�M��`۶պ�T6..N�799���O������dt�U��0-g�2U%�Fd	�:S(�$B^z|�����aл��d?    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:55+01:00" xmp:MetadataDate="2022-09-01T11:07:55+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f4e2f32c-63c1-f04c-8c9d-5c36ded8df2c" xmpMM:DocumentID="adobe:docid:photoshop:7eb11e4e-d4b9-794c-982a-5afb211b0df4" xmpMM:OriginalDocumentID="xmp.did:2ebd9bd8-fc61-3340-88b5-4d2a221384ac"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:2ebd9bd8-fc61-3340-88b5-4d2a221384ac" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f4e2f32c-63c1-f04c-8c9d-5c36ded8df2c" stEvt:when="2022-09-01T11:07:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>:��  �IDATxڕ�MKQ���Ɉժ���Ȱ��-�\TD�&
�EX��Z��}��(+�DH*تV���� �P�g�Nw����������~A����5�G�>��F��Ņ����<�g��L���&���R�T"�@UUh0���L�2�*p�����V�3 �@ӎDc`ڥ̰)�i+j�Eo�6�q0�� �����-�ZS#t��;�+���Y�X�ax�RN�^pu���23�����чc��eA8 s+@�e��j|k�f'��b���m���4L�>D��B���Z��u����H�f��ȱf���w�H%ëɵFi�.�mb����z��EE֛K�Ƞ��ꍟ ��	rJ���kd��E����m'�B�8	��~5�u~� �b��	R���o���V�15��k"���	�V���@    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:58+01:00" xmp:MetadataDate="2022-09-01T11:07:58+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8aeaf910-22e8-8f49-a756-167002efa0d2" xmpMM:DocumentID="adobe:docid:photoshop:9f90c1f6-6a76-f742-a9bc-e72d1d920575" xmpMM:OriginalDocumentID="xmp.did:7b248eee-72ec-1e4a-b34a-cac07008f40f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7b248eee-72ec-1e4a-b34a-cac07008f40f" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8aeaf910-22e8-8f49-a756-167002efa0d2" stEvt:when="2022-09-01T11:07:58+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��&  �IDATx�cd��͜���_��Cvz�� #>RcQ���_��������?�0CH6��ۃa��=pC�5���������a �����dVFbl���dpv�gE�H� g�ع��l��5`p9��o&��;���c�	�0�s�G1C���o�-��xY���F_Y���������d��V�A�VÐkK!��0zh3333l���p��/#�F�!�W<��d�۱���wQNf�� |s�L �;¶�<g6f`�`b�L�oo|�)����έuOq��v�C��g^2�h�A4���ٷ_������h+g/��`�K�.��D��� �X�K����o��������������~�>�:���~������?@�N�0y�!�3�G����?g������$�R;� ���Zirm    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:11+01:00" xmp:MetadataDate="2022-09-01T11:09:11+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:9d07ef79-553b-5d43-ab6d-5d9e4103e695" xmpMM:DocumentID="adobe:docid:photoshop:21911a6b-489e-df4e-9f01-774e35400e5b" xmpMM:OriginalDocumentID="xmp.did:f5f99420-f2b2-7f4c-a43a-1a6d24cd3bae"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:f5f99420-f2b2-7f4c-a43a-1a6d24cd3bae" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:9d07ef79-553b-5d43-ab6d-5d9e4103e695" stEvt:when="2022-09-01T11:09:11+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>>а�  \IDATxڥ��KaƟ��4���~9��d{P�P�"V�TKb!���пM���'�X-�nSG��y�yo�	�ݝz�3������}��s������l��s���][�Vb�m���^��Zg,f��,/Ɛ���A~�Ak��TR����F HW�Ѧ-�5��q,Dְ>��7`3�yG�K-y�B-J��K���Nlv�f�$�мV�O~�|��!��{��A]����(Vc��yve�|PC�"���G	L�%te��(ʪ0��d�l�zaB��t5���*����ؙ=�����X�4���J"4�0����b�C|rj\�4���+�/��� �B�    IEND�B`� 
BackgroundclWindowNameDelete in BackgroundPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:18+01:00" xmp:MetadataDate="2022-09-01T11:09:18+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d678f71f-7db1-4847-80a1-05c305c8efc7" xmpMM:DocumentID="adobe:docid:photoshop:4d358e05-7041-0a4d-a6f7-bee206a7057b" xmpMM:OriginalDocumentID="xmp.did:5d11939e-4e88-e146-a608-bae88c98b598"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5d11939e-4e88-e146-a608-bae88c98b598" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d678f71f-7db1-4847-80a1-05c305c8efc7" stEvt:when="2022-09-01T11:09:18+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>6�%�  �IDATxڕ�=,a���U?�5�+Z�DPA�t���P��b�1X-�I|��4�D|\iTz*msw��^��+�V=��}���{�
���E�8K�����DH1�@o�.;��A(J�kfJ����ކk�>!ߛ��!��rP`
�s �g������X�6G�L�.�'%�[�YYV3�F�G���z��Ŵ�iB+s�Xۅ�֔���+������t�b�W�c�7E��&to���ͷKnT�xd��<@�봣��E4XSxNX��^�ag�i�x3����t6G 40��{���X��'�'/�a𵴼�+3��%�1>!�\���K,�`���GD0���"EQ��@90��$le<�����9�6n�٘V.�P!E|�C`� b�t�}����.�X��qU���%"�H�o��yc	I�ʡ4k���潔�v�~Q�=�    IEND�B`�  Left(Top�   TPngImageListImageList120HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:35+01:00" xmp:MetadataDate="2022-09-01T10:57:35+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b6b0eab7-5227-3e4f-b344-ce0b9ec729f8" xmpMM:DocumentID="adobe:docid:photoshop:d07e584c-62e9-1746-8485-b3340c627702" xmpMM:OriginalDocumentID="xmp.did:ffde8c28-ede5-584b-82d1-a4005269b900"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ffde8c28-ede5-584b-82d1-a4005269b900" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b6b0eab7-5227-3e4f-b344-ce0b9ec729f8" stEvt:when="2022-09-01T10:57:35+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>/��@  �IDATxڵ��J�@ ����P�E)J���|
��-/�Z<��kjU(z�u)�Է�"b���P463Φ�m�
u!��~��nD$:�o�����o"aah�F�3������>*�׉0 ��V�-	!�C{�Q�	�O78w$�� V��� '"ǭ����S�0��ˣ���  �N�����;��am�ŏ����wP�F�:��7�U3L����8,�P���0��XKЫf1&�k
�Hw���R��a�6�<Bn�l���z~n W�3DmM��*��ɋj���6��s���� 
6��5�������s�m�VT(X��|���j&»_;����#5vVQ���� c�10��NG$�T��%^�D�M�Rj0Ǐs�0?.����߾w����� x1���Dn�VG'{$w�̞;�_���������    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
G  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:50+01:00" xmp:MetadataDate="2022-09-01T11:07:50+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:861cdb4d-c261-6245-b6c7-bb3f3ad7f4f0" xmpMM:DocumentID="adobe:docid:photoshop:bab765bc-e4a8-264e-bb48-0f973dcd85cb" xmpMM:OriginalDocumentID="xmp.did:852956c0-5101-6e4b-9e6b-f9cf5676a668"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:852956c0-5101-6e4b-9e6b-f9cf5676a668" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:861cdb4d-c261-6245-b6c7-bb3f3ad7f4f0" stEvt:when="2022-09-01T11:07:50+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>I���   $IDATx�cd�2`5p��Aj�J̠��T�򨁣��@ ���H�    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
�	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:22+01:00" xmp:MetadataDate="2022-09-01T11:07:22+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:6f7bab71-321e-8d47-a8b6-7d95717caf93" xmpMM:DocumentID="adobe:docid:photoshop:4bc883b5-3d72-da4a-9ceb-c582b08524df" xmpMM:OriginalDocumentID="xmp.did:e7087dc5-2d05-9743-b387-699857a51088"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e7087dc5-2d05-9743-b387-699857a51088" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:6f7bab71-321e-8d47-a8b6-7d95717caf93" stEvt:when="2022-09-01T11:07:22+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  yIDATxڍ�[hU����mg6��]����������"
y��Z
m�`�}����`%ڗ
�Z����R(J�T�,i��4&��d���3�x�m�!�\����}��������/QU=&��qBPW�ƾ�F���$��I�g��J�f#I�A5(%*���*�	��ޱWw����i���4oe"q#�Rp�"�R�/d��Y��*��JW=(	����/k���Hԇ�Ҝ�����M'�`�p�lg��I���/��y�Ŋփ��cx�c;��2�\�gW�J���~���ܗ��M��Rj�L9��lCZW�ƕIMσ��ˆ
����,&Z�D8������{�8ښą\�u��g< |�b��Jm �\�9�ւ���>ю@�{�b��^u�|�9/~D٨���bl�� ��Sg�������b�k�S������e��-��
��w=j���,zRF]_O����Ȱgh����O!圆U��Eز�X��Ο���<eM��t�
�ߕEw�����M��[L�"��>D��an��jR�"�8C���	����>�y��Ss�I�<���%��̸x����&�}��\h��kT{-��:J���+;E�y-��U�����ǹ)s���]dBC�R��*X�S�ca����ڽ����Y1�hh���p �[�#�9jT�A����O�Q�Ț��ۀ*�	x� ���<h?�H?Ϊ�V�%֖_�S�bOj6���>,T茮WX'����D��Ak�P������ixs�z�Y<�A"g�������K?��^2���X5�D���}�*g"��q��>��a���3�_>���㖁a<{2!���G�'IPaK�����N�D�Rz�_    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
�	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:25+01:00" xmp:MetadataDate="2022-09-01T11:07:25+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a1fffd4d-344c-1b4e-83b7-02146929b990" xmpMM:DocumentID="adobe:docid:photoshop:120196e3-c93c-5449-8857-5af7709771e2" xmpMM:OriginalDocumentID="xmp.did:5a02b2b7-9209-234c-b44c-217623602898"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5a02b2b7-9209-234c-b44c-217623602898" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a1fffd4d-344c-1b4e-83b7-02146929b990" stEvt:when="2022-09-01T11:07:25+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�&y�  ~IDATxڝ�_h[Uǿ������Ԥ�I�i5�,�aCP�|�)>�>�E�����@q�EE�@Й�(Cج��UiZ���צY7g������='[뺦�x��;�w���߿��p�ؿ��3�>Na����� ǡ
Νp-�u��t���ni���T���x�$<aq� p��m:����Ys-w޵���O�L}�O�䕍���:�LR{\��R�Y�Q55zKv-(���ܺ�7%*o��kÞ�qV�q�f�}V�>���}�gd�1Y�?�'�Z��1?���J{O�A/�u�v��m�j0sxj�w�gPR��0/����S�I��(b��,ÁQ�F�=��:+��d	���/��S=a������|��c�f�g�d#���_�pF!�`)��#w�aSݮ�*�j��=���َ:t'���Ϧ*�no����#����|�-ޕ�@؋C3�x���e�C�հ:[�b���{}	F��|Q���6�|��C�3�i=�W���ԝ1u({o�,���<
K����C��ÿ��R���������]}u��,�"�#�����q�7�>#����%�~8��[)�ǿ�x�t�m��?�m�G�o�<����F1���E�Eb��Ņ���/E$y�/�#���x �4\��dnn*LⅣ��7�C�.��F�av���������R���Z��y#���^��ʈ�Xhc�qsk��1^~�}�t(RT/��=�9��9�=0i�ĭ��n�sp�]?�8nµ����Ͻ���r��P�9�VJ��ц��6�,fO���B�����6Ls�nt����ni���.�Lf��|���m �_�[7��t*��U�V�i��.�/��\( ��}|���� x��i�ze	v��"OX-c�?����{U�`    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
$
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:31+01:00" xmp:MetadataDate="2022-09-01T11:07:31+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:51f68140-76f7-c04e-ae9b-4331960aab30" xmpMM:DocumentID="adobe:docid:photoshop:02e3f29e-a481-c647-a132-1a4222b5d70c" xmpMM:OriginalDocumentID="xmp.did:52b5723f-8145-4d40-8f90-f3f521782e7e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:52b5723f-8145-4d40-8f90-f3f521782e7e" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:51f68140-76f7-c04e-ae9b-4331960aab30" stEvt:when="2022-09-01T11:07:31+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>vX  IDATxڍ�	Le���͞��]�h�E�hi�BUڈ�Z�#I�V�����xT���D��Z�F��D��4hӃ ���+JZ97���2�����7T�
4�L��;������}�k{�gB��D�+SU5MUaeL�Q/��򁧧�k�G����'����ꘓ��Ę��P���!�iZ�0�R%�O�ļ�G3����;����4Y�V���FU�4UP/LI�8��)��A�	I[.q��UF�Ⰷ�m�����e��;<]5)]����u���~j��B��EX���p��Q��a"��JIo�m��&T�6�,7e8vA���rb}<":<yыơ)H��/5z��޵�g��l� ��i�=7E�4Ύ�Q?�~�]Sd@�=[S�Ϊ�d{G�ś���tB�s��<���k/+����?k�YV�m��kMz;�^��Q�����1l��)�Ki���ÌY:���d98t�E|��ṛ#18#��n��(htamgL���Y�'ԩ��rv��T�HUH���x?5i��s'�l��?y$w_������i8r���EA�b�̗J���Q�ٔ����-��.Ao&�~8�n%�Q�#~<�|�F6�}��r��>6��]��`��_��w�l��/��;EO�z�ު32��l���� �q��m���4�vDl~c/��7����0�b�-�ߩ�����C��]��,N�D�f6D+#�05�����B��|�{ �aX�a��ib���]���5��u��ڀ�;(i*��z��|�5�%���/�t�i:�@�G��_�D�#�2��ǅsw:$K���Hf������k�����[�8��g��.��.�n�$i�%4���Sw@�}�*o���,�e��9|C��J�7+�<��f��R�ѓ!F���x9DO�؊vC�\�/�7�g���.	�YC�n���6�繰�2�('��];���ut@�w���KjV��81�N�=*l�_��𝨈��ѫ���@�&C��    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
�	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:28+01:00" xmp:MetadataDate="2022-09-01T11:07:28+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:47bc6c71-0dc2-3f48-8f21-f588a06d881d" xmpMM:DocumentID="adobe:docid:photoshop:dbf92cce-85ae-4c45-aab8-e1ac7899fd04" xmpMM:OriginalDocumentID="xmp.did:c261ee3e-fe3f-8448-8ae0-d3d5900bdc35"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c261ee3e-fe3f-8448-8ae0-d3d5900bdc35" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:47bc6c71-0dc2-3f48-8f21-f588a06d881d" stEvt:when="2022-09-01T11:07:28+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  �IDATxڕ�]LW���������
���"$j)�Mx�����Q_4*�T}�Ml�4���4Z%&�(mb*~�VC�������L�ݶjAfW�ٙ{{g�[)�œI�=w������l���`��uT��s�k8�����.n�������
#/&����$�˒������BA(��a0�1�G3In�7����8P'�3\^�+S0��=�|��1�4-c4��]�'�����uw��J��V_�C�����u�Э^����|�'��[kE:�)W&��,�`��Y�<Æ�(�ÙT�b�o�� }�V0�U�T��0�P��w(q���G��$L��H�m���w�G|���0��3���E��Ha��X�� C���.� 6w[E!����]�%����!�L?��ҺŴ����~��v��8ZӢ2;$l	�14���%�XZ�FS���y��11�O���5t����.�C�P[��?e�L|{+g��1������������dȦG	�,��BӴhNe��6��T[�o��P3͝۱�3��t�{aX'@�,|�c9��ŃD-���V,)�[3��{�yV��8=r��T<8�x6����cl���v	%Ʋ�,����up)r�?x�:�jO2�X��Mqа����
�.B��ԋ�?t<��Z���W��kk����9���Ӹ�?2�.Kh���Jn��n#�1m��[�'�q@Ut@��9��+����K�d\�?P����pP�u�i�/߽���Ǖ�wDbh���I0�[Qz��~���W# �������)�����m1-|����u�,_V�4�hJ@��ͫZ�3R�ɮ�0kz!�Oq���l���A_���)m��+�"ӽ�U d�肘X��1p ��옿
��Lf5�l    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
$
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:34+01:00" xmp:MetadataDate="2022-09-01T11:07:34+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:39076e47-50ad-9744-b953-e0caea6e9324" xmpMM:DocumentID="adobe:docid:photoshop:69ef7004-ceb9-704b-9e15-039c68d19f6b" xmpMM:OriginalDocumentID="xmp.did:f9f27a3b-28a3-074e-babc-9fbc89a2f251"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:f9f27a3b-28a3-074e-babc-9fbc89a2f251" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:39076e47-50ad-9744-b953-e0caea6e9324" stEvt:when="2022-09-01T11:07:34+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  IDATxڭ�mLSg����޶�ޅn1���Y�{���*�����4fn��,����A�鶌�/�֥�ut �i@�6d�&ns�f����mo{[z�^h�}�ܜ����9���P� �^
R5Ñ���R�0�ĳ���c��d�t���]�ږ�'��YӁ��t�ё1V��V�K?D����f���E�G�����[7M�MM�w���Ne�w̅�4M��i?��π���}� ��8��8��Gػ���z�mk>�1���3_��ϕo��<R�W;?/����
J����	%UN��}����)@Ú���_X�B�@Iz��x�N�T��Y�!��W΁=Y���ŏɞ4�t�V��KKW�ݚ��rR��Ė}f��m#�����΅��jH�b)������~9�@U�Y�F����?�����!����L���f����vj��Ga��b�v%h�FpPpn�� ��a������Y��}�[ׅ�}�T��z�����V|6mނ���P�T"8;+s<Kr�;�9Xk)�S��-�W6�}"0[���-�˺�H'y�>r�������t�S�{g5��E�؟?�Y�'��]ގ�������"0K��׺��V\�H�|+Piă�.]FY����b{�6Ȥ�q��X�C2 �<�W>�=	$�۹�X��Л$  _�zp1ٓ�0�a��j�9PJ"[Ձ��]W�?/ِW`1ט��@���$��W}g����r�C� Y�Ol@]���8<є����s�4}V����R*Μ[�	\DJ���8U�g��}[���n���7u-G�O�{u��.S�q�.��� O|n��pJ��������a{�����W�f�ݛ�yK5/y~8�)C=a�������'�r3�^h9(��&��|&55�
]��;3hwvv
�l6�z�n__Q�VF��h�ZF�� ::J������mmd�xzF����]_�KZF���P�H<O�|�8q�ʤ�$דn�kks��.�{)��}��Z~    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:56+01:00" xmp:MetadataDate="2022-09-01T11:07:56+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:026a5789-985f-5d47-8ae5-3c152a2c3138" xmpMM:DocumentID="adobe:docid:photoshop:5bb8c5f8-e193-3a4f-a9e7-9ea29d189eae" xmpMM:OriginalDocumentID="xmp.did:7850f5eb-cfc1-6b4b-86b9-02544801f4a4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7850f5eb-cfc1-6b4b-86b9-02544801f4a4" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:026a5789-985f-5d47-8ae5-3c152a2c3138" stEvt:when="2022-09-01T11:07:56+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��ŧ  jIDATxڥ��k�Pǿ/���8ש�tʮ
"�ŉ�n�����a���@��<���!e��M���AD'��m2
-��[�i�6i�_�5v�ͪ{�C�/�����G�ɸ70d8�uV<���|[� � �:���!�j^�Z��-�.�`,������(��EL`IM\�	e�NF�˅�g��wOÆZ����3Ќ�2�h�m-��F�y�7n%��>�9tr�z�]�+E�?<�H�S$�YY�+Mx�𚷁�qJ#~�O�!'�툊���G��w�Q{P��/5�B&��q��#8J}�#+�i��{�3�HG%�j͡A�+�6�F٘7[�~��E~��[� S�d�x�&w8���]�IBW�QS��l��w	��p��� ��q:���ǐ<�e�����s��.q3��D�[X�Z���ŗA�D�!��c*��	���X����K�	������4��U�����z���~'þ�m�ƽ/�Yj�i*ʧY{���|W�7rJ��"�^���/��� {P���4�.͑́yN2�}6ڽ�8��ww�d��@�%�T���c���t�����7����}�f�Z2    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:59+01:00" xmp:MetadataDate="2022-09-01T11:07:59+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:83d6dade-5656-8a42-a3ba-9cd23c35b21c" xmpMM:DocumentID="adobe:docid:photoshop:6943318e-c4f0-3449-a1b7-cc92fb7f8bba" xmpMM:OriginalDocumentID="xmp.did:d3b85b71-ce7b-2b4c-a61f-971d9a9df163"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d3b85b71-ce7b-2b4c-a61f-971d9a9df163" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:83d6dade-5656-8a42-a3ba-9cd23c35b21c" stEvt:when="2022-09-01T11:07:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  kIDATxڥ�OHQǿof����U'�-��С�'�
�"H�K�#f(��kD7oH�!(�)�.aւX��f$$���ݝUgwgg�ݙ}�讚��<�o����=�#(S��!Z�mZM�nWǧ���V��������q��1��<���Ο��HpJ
��	!�t�m/b���۝7���RFn�Ǚ��������� ��ߎaEܜ�ۮ�5"˲h�qm��~#�j�+kx�*�h������Rj�D�툗'1�r"�3��u�:(8�V�ମ ����-��8;#�EWk�|pT� ,ar�Z��&�:F#%�ו�7SEn��s1���lK���Eن�%���k�a�T�� �-voφ�C/X��*V��(�@[����k��dx��M=��AuC�eG�X � �á�O�-k�Lg��d
sF�59�:�@]1R�$/o��׿u-I�%�,���zh5T��\7����1T)	�JU�p<��?Y�{Τ�$GQC3k=t�'�h��0�4W��&�ӚNO!Т����[{������ґ�@ݠh���E ���VgzJNOk�X�_
B�G�Œw9i���##
�Fj43����>����2N(b�`v�h�X:Y    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:12+01:00" xmp:MetadataDate="2022-09-01T11:09:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d388fd30-6b31-064d-b3d2-82eb6f97625b" xmpMM:DocumentID="adobe:docid:photoshop:806bf7ad-fc45-8646-bceb-ce24e6f2af7a" xmpMM:OriginalDocumentID="xmp.did:50801632-0a6b-a840-8b87-4bf6c0099d55"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:50801632-0a6b-a840-8b87-4bf6c0099d55" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d388fd30-6b31-064d-b3d2-82eb6f97625b" stEvt:when="2022-09-01T11:09:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>]sS  �IDATxڭ��+a��ow��h�U�)��(�QԺ�{^b/"�6ܔ\�$�����=n�7EyY/�,�v^3+/ˌ5򭩙�7���4�c������ߪ�:���w�{���j�s���E��5��Vaw��5js��C4�0��}���m�sC��*Hjh��G�k��B��k�-#�Z�\K5l���L���I��-���T䵁@��6���i��P.A�c;l!
�e�4l]w�z5�-�B�$	w��cX[>��-�Ns?G� �g6���G�{��b��7T�SE|=����z!w$��`��yP�~jG*' +X���QjZJy��m��JQH
��y"�{m�C������R�6.��L/���"ri�7�E�H�Sb>��yPo'hK�xɲ 5�A·��q1|�H�C�k_�h|g�n?�n�|�fs����    IEND�B`� 
BackgroundclWindowNameDelete in BackgroundPngImage.Data
  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:19+01:00" xmp:MetadataDate="2022-09-01T11:09:19+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:0b77d393-b5d5-a540-9862-7c16c9604ce5" xmpMM:DocumentID="adobe:docid:photoshop:7323815a-e372-0e4c-ac3a-b14b03087c93" xmpMM:OriginalDocumentID="xmp.did:a7567725-d612-374e-8978-f22fa6a4e34c"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:a7567725-d612-374e-8978-f22fa6a4e34c" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:0b77d393-b5d5-a540-9862-7c16c9604ce5" stEvt:when="2022-09-01T11:09:19+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�ކ  �IDATx�cd  ��>���_ƿ�,,L���1�X_��ًW���0���	3�b�U�n�{ 7���gddd��"�d B�Ꮵ�+V񹈕��AI^����C��Ԉ�dA^�s������0ׂ$׋LL���ژ.�ċ8]H���a�cDz�d����i�����r���P\���	�]E������Btמ��b�������%����A�ݯ�e�c�������Ļp�2�y�r��^�g��I	P�G��0|{�ʆh����0ܯ�a������_��_?��Uyr�ݛo�~8]�s�xB��E�����O�x���/�a`��B0�{��aN��$={���wl���f6���dxE�=��$c���D/#�_�)In�Ͽ� ���,@c$P"����T�w��~�����_��^�g�b��ƺA��E������0�_�����m����a�� �PVf��??~� ��a����n    IEND�B`�  Left� Top�   TPngImageListImageList144HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
b  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:36+01:00" xmp:MetadataDate="2022-09-01T10:57:36+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:476080b3-62e3-864e-915a-47b66c957534" xmpMM:DocumentID="adobe:docid:photoshop:182e7d80-cad1-214c-a9e1-1b656de377c2" xmpMM:OriginalDocumentID="xmp.did:581990f0-e9f9-2844-b56d-bd917ec672b0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:581990f0-e9f9-2844-b56d-bd917ec672b0" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:476080b3-62e3-864e-915a-47b66c957534" stEvt:when="2022-09-01T10:57:36+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>dn  ?IDATxڽ��n�@�g�4���5=�V	��|@=aY�U�3�7��"������Gh8s�*��N�m��ìc�6n�(�e���3�k��0͇�7c~�Y� �{��W+���ޮ� ��w���V�M�tޮi�4����N�5꒒�`� y����C����)�h�:u�n�d�8��ヽ3#/x�����xb49��#%7����9��~��P��T�J�a�
-�����<�~�P!H�*e�b4��%&����]�7���G�6J� �J&�f��t��&@�����
RI��k(Qa�!���a��8z.%HS�h��+���K2H�m��$x4|rA�s��$Pla���c��@���:d�q�Dq�E��������#������DE�u]�����1���r�t<���zW���SM��d��*�DQ�-��[x���R���+��e'�J��J�
j	�V�����G��߶k�	�!�J�s�I)HWB��>��s��%af��eYxVR)U��j ���pD�>_4fgػ���B���V�yr�?��z�.�jȌ�ENA    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
K  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:50+01:00" xmp:MetadataDate="2022-09-01T11:07:50+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:375ecdd0-9fca-6e44-8e6f-e5190740fc98" xmpMM:DocumentID="adobe:docid:photoshop:48e9df4f-c528-184d-bb90-8e84a567edf0" xmpMM:OriginalDocumentID="xmp.did:86b9b7b2-08b0-9f4d-ad35-1e46758e57e4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:86b9b7b2-08b0-9f4d-ad35-1e46758e57e4" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:375ecdd0-9fca-6e44-8e6f-e5190740fc98" stEvt:when="2022-09-01T11:07:50+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>� �   (IDATx�cd�1`�`ԂQƂ��4sxZ@U0j��� �uv�&    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
c
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:23+01:00" xmp:MetadataDate="2022-09-01T11:07:23+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:76554e46-2940-6446-8c5d-41201dc69565" xmpMM:DocumentID="adobe:docid:photoshop:7982d76b-2c09-c24b-9d96-a9fe01b2a6ae" xmpMM:OriginalDocumentID="xmp.did:07a46818-2a37-8342-b693-390c66bb8de5"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:07a46818-2a37-8342-b693-390c66bb8de5" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:76554e46-2940-6446-8c5d-41201dc69565" stEvt:when="2022-09-01T11:07:23+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>c��  @IDATxڕV[hU�Ιٙ�d/�ͮ�Msi�F!	,�
y���⃗Ҥ�"�Uh�<��̓ZD�6
!��*���`�"���D+�l��b��^�;{�3�3���ɦ�v~���|�=;��`��.��w�P�
��!<�!�xW<�=�G�B�.���%D�pʪ�q8%�@�eMi��l�%�4;j���"��|�P<�.wj�B��s�/땵�1��M��PK}[^�]��2��ViN��\�\<4J��)]��6~�%��s��?�Y�n���eh�p�o��HE���H�b����1ŭ�r��έ��p���>����u�cF�e�������{/�49�4'����B�*㇙8��6aۘ�G6a�4��IP��@�[�y��o8Z�SU~$���G�O2k�1�-�FF[|�S�=�|5�^�T���J(��f�12��N�Ef�I[F�p�4y�x��t^]@�x�io(���B\ѳ�'��Z�<�WP��	���~f��w!�	^�\[!���Իe���"�tk�6�5<��xg����}Wqaz%��A�g�*K@q�i�E@��E���)2m�Ʈ�V�ȡ9N9�N���۶a_��M0�E��"^��Ӈ�E�Vb��`)�k��;u���$�͌Y�{<2�4EœZP�P�س�V'HJ�HtQ�=熡���W6�%8�k��%L��Ǿ���aOrՇ���|��͚m�	N޹��{���3��/Q�hC�!n~8�|e�F�\����/�BNx�HK�<"=�CٵcV������t&B�OH?��MŝD(�8$��$V�ĉ��ݸ�!j4p��E�cCrl�%����kE�x���4x�a����/rف�ɞ3�hq#�l� 78þ��&l&{���wU���E���+:+��)���"8�; i���:V���!Yg)~$/1�to�?����jФ�O�	��Hc��-��G dכ�ZI�/j�̭�F�����S3R�e���NĆ�&�d�;��T�{��K� +�5�c�RK:AzAJ�i�p�<�lt�:sC+�z��{Br�i�H#�g���߹��;��x�m�/~����e͵    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
�
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:26+01:00" xmp:MetadataDate="2022-09-01T11:07:26+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:51edf77f-337d-df4c-9412-c02490953f86" xmpMM:DocumentID="adobe:docid:photoshop:38f42b90-13ae-6648-ac1e-ffa02882af0e" xmpMM:OriginalDocumentID="xmp.did:c0055a1b-163f-6548-addc-8e97eea98b83"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c0055a1b-163f-6548-addc-8e97eea98b83" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:51edf77f-337d-df4c-9412-c02490953f86" stEvt:when="2022-09-01T11:07:26+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  _IDATxڥUmL[U~Ϲ����Җ~�BA�:u.�3��_��g�%����h6�1�?�_��D���0YLH�E3��e$n�"�l�������s/�QC�UϏ6�y��y��� ����_(+s��F��ã���k�ম�é��P���<�A[�����B��²���TYE�@Jʂ*h�j�|g�O%Gg�GN�O1@�A���M[�4�bF��|GC��_}	[𐳎猈����R$�L8�!���W��%0jnw�5��X��'OT�^_�<y��
����d<V]�'�D�:cg��*Y�x���l�2����m��e@\SU�ߞ�l�/H����%�ߺ��pAp0��t�Y�z/ǯ,�>��CN+�s�-	�����Z�i�~;p� ���Z�U��'�`Y���h�'����FW��̨� ��Ws���C��fB�Ѽ>�IU#%��f`����88��q?-���	���V�ngdh'�ˊ�72P�J���ӗy/����p�����3���ٔ�������N��I#$}�Lz�T�)�y���Мq��X���3�j`�0������+2���p�� \����nAS�w�Nm�hf�����d��uP�Y�}�S��^�.BR�N�!�}��,���9
-�(�f߻p��D2�������V��qS�u?L�4��w3��m�#��]/���{��ܪY�����`W%�kwT���i�w�O�[遚 Q�\,*e���.��ڋ:au2<������'!�y��t���'$~��,�ݭS��&xu�ӽ�w"w��M�NB�04ES2J��O�N�GSt��l��o}�g���8<KkQQR�:\]�p�,*&xn�m=�� �C�=x�lM���{��#�DlШ�1c	Ul�HT�z=���R:*K���%(�7ӟ���Q��c#AL&ůڦ�yc�_�'��+5��au��b�U�Z�W�Q%�v�N��p��ƽ����2ܵ��x��#GR2�&���rG�j�̈�!���c��K"0�<�u"w$�Gɚ�+ǆ?�s"Ox�_�x3s��B���K��O!�t�i�K"8�?˜E*|��V��#ˢ���Ϗ�5^    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:32+01:00" xmp:MetadataDate="2022-09-01T11:07:32+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b0e45b43-f18b-2d40-a2a0-54ec0206ab48" xmpMM:DocumentID="adobe:docid:photoshop:20f8234f-b20b-4843-bcce-ed633a0eda9e" xmpMM:OriginalDocumentID="xmp.did:52bd6386-6c2a-ce4c-a84f-7df669a07cac"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:52bd6386-6c2a-ce4c-a84f-7df669a07cac" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b0e45b43-f18b-2d40-a2a0-54ec0206ab48" stEvt:when="2022-09-01T11:07:32+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�y�I  iIDATxڕ�kLSg��紧��B/P��:/�
��2j�%N�6qn¢q*���%ۗ��9����͈���$���p\4YD��"�(m���s��Ԩҽڼ�m������y)<�bJ�#"4��MeC�$Q��%�B�ȋ']�����.����7���(JVʨ�J��ae

>  ��w<�G����Z�gT�/@©�m��H#��4 �E@|��x�����"�o,+��ğlZN��2��cC�d\$M�E�q�y��|�%'��Q!�#uQ]��f4�C��$�CfL>����~�߀�a7���x��"R�;"NɎf<#*���IZy���n��> n�d'���x���0&�a��+@�9f�r���¦�.�'���L�5" ��١��iBڿ�8`C���Q��"޺t=�79�w�St#KT���8z$�&V���&@A��ڇ���g��s��H6j�&V� ]�b��:m8�a�����^�{� ���oT!��,&ܿ��I�T���k����J�=�j���ir%��8-�L���۬hw�p �(���w�V[�*6���QKa�@N|�yx�A���]A�)|�������F3l���ɱXbPKF�x*���Q}_�d���#&~<T�>�"e>����*8�}����Z�.���f6��ph������QR�N%��a��$vQur��E�������F��
xkd�F(�̆H��ߕ��?kx���v�/I�d��4��\���6%R�>-K��ك���=�I���"ġA؊VApڡ�-��`>(�џ� ���a�\t�u{��r�̢��B��6��(8J)�j"� ѷ��cdZa�+;?�/��q윷��;۾�p_>f�T����Y��#P��4%3���R#cd,�����=�L���t�Z�lx.�%��#���Х3�l���<֌�U����;@=_�O��y�L���l�L:qr�*����C�=,EԦ��/ZK ����o�Ղpw��|� /ZuiJ�٬֎;҈`�m�f^}ћKѿg\u� C�Y0�I�dO�}kp ,��tem�X.ô� ��,)���6�B��c�~K ��`�&�x�*�U��u.�.�rX�����>�Ҍ$�aox�C�r�����o�ZIöJR�q�Z?�����A�	@Z�^��l�������-�drx���)\�B�|=;��W}^txE����a�(Ra�ъ�(-��N�Dk�/ ��h�C�`/�G{���`����3�6 �j�O1���"9Z���J����.�8D�~���F;�ܭ"\�^OU�'��dh��G��2H�-�(�i�����i�/����    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
�
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:29+01:00" xmp:MetadataDate="2022-09-01T11:07:29+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ab0d6e3c-bcce-9f44-a750-4581f725a497" xmpMM:DocumentID="adobe:docid:photoshop:05cf6a39-0539-ce45-a23e-86c81e1119ba" xmpMM:OriginalDocumentID="xmp.did:529115d0-c3dd-3744-a1dc-1e55436072e9"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:529115d0-c3dd-3744-a1dc-1e55436072e9" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ab0d6e3c-bcce-9f44-a750-4581f725a497" stEvt:when="2022-09-01T11:07:29+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>ʥR  ~IDATxڕU{LSg�}���^��
����1̀���M�Zs��\��eht�ef`�`f,Q�&3�x�973�D�^����@�% Aǣ���Ƿ�^���z���;��w��<.�CY�j�O8R�dJ��:;�i���d�Di�,���P߱�]�>$�h4�y���AH^��݊�B.�/z��GHl�z�p8�:(�����Y�*pOx\���´�� �l{� ��lx5b�)�8�,�Ĝ�������Պ *�a�;���J���O�[���P�mğ�ݘ��L;�&�V�	aї���1F~%�[,�8��F{��!tN����ܲH���U�X������9���pu��� \�š[w4���!>�Z���$6tN�����rΡ ��(�Z��)����]���Q��;#N9����ST�%�'
�?�q��n����}5}�}��q�
�H�baq��A���{�Ѩ�u������Xl���K�6�(ʐm?C�	:�8��<®���=���� ���.D3��vǬ±�H�P�{}��Έ��Z��K���J�t:��IQ7c�����Q�~�Tw:���.��J~��W�)Q�mҜ>���8�0�����2�S����&���B�gujfg/���/�Uz�)�7S���U�G�H���m�*�` 1� .U^s/FO�:6���s�)�z+oD��-�(=~�����g���,�/:�9=�	���6��룰=֌n����k�/|�l�,ٌ��l�ɚ|����Rv,B'��*X$���������ʐjN�vw,ap�b1�A�5���$��3�d�{�m�v���^���D��!I��ŏ\>�i����΃���;J���= d��q�5M��=V���nG��D]ɱ+h��! k�S���h�K���.�G���	��c��\c���@k0��"������?@r>״��H�3x� �G�ѹ|�Ъn�]0�X�XiK��nI©�[}���O}8��wlO)�޿z2�՚j2�MeE=�V��C�<��\��S�:��$K^dt�J||J�ހo��u=�������!J���6ы��=��;��@WbRꋬo��g11l&�E;%JC��~	K��?M�9"Ϡ�>    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:35+01:00" xmp:MetadataDate="2022-09-01T11:07:35+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d20ca985-7583-4f49-9cca-3184c386e1fa" xmpMM:DocumentID="adobe:docid:photoshop:b92fd3a9-7f78-0048-b0b5-e11bfed08904" xmpMM:OriginalDocumentID="xmp.did:7751f063-a01e-ac48-a206-5b0fb2241355"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7751f063-a01e-ac48-a206-5b0fb2241355" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d20ca985-7583-4f49-9cca-3184c386e1fa" stEvt:when="2022-09-01T11:07:35+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>.���  eIDATxڵ�{LSwǿ} i��3�L�)P5���FEZl�ن(��[�Cd�f���-�E@&\|��n�Z��m�TJiKK�{w�-T���_��_�=������w�a�$�W9X4��bM�1<<��ʎ���C�D�^oҖ����l��jPU6�Q���r�D������_�	��p�9�E!_�����B''��<��CG�]��r�uE�@���C�t/DDD�Ne���7nH�sXa�o��~�q�H�	l;gp��`=s9z���GK�ZZo��W�/��=��\@xd��Ͼ5)1A���7A�(�Ӂ4 ����o^lWlA��FSىr�V�54�u�в�7'���j	W{.Ʈ6�3�0`}g����_W�3W���S�=g�r=�\�ٜ9���ڞe�X����b�,���
��-�e�?�WH�o�@٘!W?6K�{��������Uy�X,v�;�t~s��IZ��~��,��C��l��/��5�L��N=`�s��փШ��l�ux:2�lժ�{<�`yd�ڹsC��J��Ϯ�4נ[�F���������¨K�2CFr��7ܦ E)�3!Y|�
�O�^�����@LBR��i�Kxk`���1f9�p�3ٹy�Q�<u�DKVb�E�Uс��� Ês�� />
��%�~��8���O�:�e��{�1��C�d��\��f��[�������۲3����8�!�2��'�$Hp��P%�E���G5U'�@Tt�����x���'-�!1� �-�q��K�В���2����=~:�Y��
'��i�g��<����g��6@��E@��X�8-�EEe�\.�rs���m9Sw?Y@MH�B��ͩ��c 1q�]�{�xLӗ��+c{m�Q(�9fHww7�����gZ� m~23��Z�����c�S�b���RS����������d��N��G�+F����p�];a����P���]����B%I�Z���#���4��Ӷи�Cg���[.BW�.�',J>�}?���F�hV<��L�9�<(��m?�#�M�)
Bb��-h��<��iI<����f��)�_��?ߡ�{<ŒhL���f�B�s�f���������-����HGȊ�&)X�*p�h��V{{A��:w\���?�U�#Y!�,޸ݎ-������O������*{����r��Mj���8EE��N����K�d�i�J��OX�-m��l�}}fx�MJ�uqv��1���n�U�Cܹ�@�X�3�ez�l�ف�f�5��`S�����6i���A�B�@����2�������o�O!"�`08Q��Vt�g��5j�q�v��M�U�xtv����    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:57+01:00" xmp:MetadataDate="2022-09-01T11:07:57+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:18df26a9-5323-444e-99cc-a6e27518d450" xmpMM:DocumentID="adobe:docid:photoshop:5e72ac25-e678-2943-b486-3117fc7b0bc2" xmpMM:OriginalDocumentID="xmp.did:c636900f-777f-2045-8d5f-e5a13c2ce88f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c636900f-777f-2045-8d5f-e5a13c2ce88f" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:18df26a9-5323-444e-99cc-a6e27518d450" stEvt:when="2022-09-01T11:07:57+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>j��  �IDATxڭ�_HSQǿ��[�|�$H�%��(� 0�z�z
)C�!|������$��J��E8i	.�(�qn�ͻ��{����6�v���r���~�����s	t�ݮ�#E�\j�{��HV8�L����`4C��M��p��
��)�������)�I,����paH���Δ��mmV+�DɆ�s4 �g ���~�R,ۏ;�/@��CoFVt� ���9a@ӹ�T@>��5��x��&+ocz����$s�q�a����ƍ�]� |���x�
N�]椵�3o�f{�	�Q �"*E���8����:"4�}�z��Dκ]^�w`�03�b��8' 8Mfs:�GMO9,e"$��'���dO���\�(����G\ $���ێ�*�� 2�R���M�*D�l�Hv�qv��\�s�� @��c�p-Zr�����8�50��b�9�.�a*�oNbk\<�[�$��v4�gb#���w���K�" !/	���8�*�����ᱻ���o�4� �
�tq���C��?�T�S�YtY@���fߓ�gu9���f�a��D3�!�'�)CPVP5��]��A�Mkp e�Bt98�]����
��-�/*k����^��
�;x%�L ����q�ނy��h�)k'�U�/i��ɂE;H��#�y���*����_ ��#��F���_��0�	0�%nF�iU܎V�b�����RVW0@    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:59+01:00" xmp:MetadataDate="2022-09-01T11:07:59+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:2599e910-86e2-4f43-a036-737f19759ea8" xmpMM:DocumentID="adobe:docid:photoshop:bba4275b-a819-614b-8e64-863216c5d3d9" xmpMM:OriginalDocumentID="xmp.did:d39576d9-e813-5a49-8574-ca8b2d2c0334"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d39576d9-e813-5a49-8574-ca8b2d2c0334" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:2599e910-86e2-4f43-a036-737f19759ea8" stEvt:when="2022-09-01T11:07:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��'�  �IDATxڭ��KSaǿ�e�չ�M�vӍ��7&Q��!袛^!î������
2����H)Lщ��N�E���2�9�Խ���3O�(g͹�����yy~|?���<�2���N�@KJh�knj��������y�;��A�t$�q�2!�
h8}}�� �
�}� D>��`A������" ���M����B�ը�8Z_��RK�@� ���B��%G������t��F��=�.�Gk�kܞ�V;�۽��k%���[�Wh���0�G0��RI���,����y=>�'H(���ҐP�Hi�{�J��bEqp�x<� R��z?��T)���U� 	�@�YXV�:��5�Mr��yϰj����|��E�c��rWA�U֟���PRe��}Y��D�eK[9�v��YdD�͜�u&�k�G��lؑ���~/b�!#h�!�����ζmw��5���$���{@)�4d썛c�q[n�N��/�բ��[��B��ca�z�D�k���p��2�:�l=>3~&��W�3f.��2�;��$�sEvt$Mbn�?m�-��@���_�UH��9�\Lje2��3�j�����e�FPT��Np5�_{��_��VX*�J�3��Tp�I�K�"$5~��m��)�����P\Q,�o,��,.��y���?>6^�k*�p���%��X�'�]���k���o�\���#.�_�q�owF�;    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:13+01:00" xmp:MetadataDate="2022-09-01T11:09:13+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:988796c7-bb9a-8d49-ade5-79e46755cf89" xmpMM:DocumentID="adobe:docid:photoshop:74db8562-b0ea-1240-b5aa-5bc16e547f68" xmpMM:OriginalDocumentID="xmp.did:fa44911e-0a74-e647-a444-9abc7aa41c67"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:fa44911e-0a74-e647-a444-9abc7aa41c67" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:988796c7-bb9a-8d49-ade5-79e46755cf89" stEvt:when="2022-09-01T11:09:13+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>(�~  �IDATx�c���?-#�,�>k)6�*��NO>B�)��D�>g�b6V֯?�� d	��z{0�ܵ��%d[ R���k��`� d . R� YB����Y��,T�.K�0R�[���|D��݋g��mgd�"胸������ƿ����	�"��l�/�$�ڀ܆��ǀ YB��ψ20 ���+p0�+�1�s�a�A�Q�� ���KB�)�b#��{�z�%�L�(���2��@�I0�j�!v)�h�v���!,8����?�|pT�b0�%Z��.�K�s2�}�?�>��d�|�x\�j�P��?����1+7�sp�#�G�Q���������mt��8j?$��⃄�"��8�Qig����Ȉ���"(�fBW�T�P�jvf�T����H�2+�]��S�A�M�OY50"vC}������k���2�^u����8��Z�v����O>(��@  ������l_    IEND�B`� 
BackgroundclWindowNameDelete in BackgroundPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:20+01:00" xmp:MetadataDate="2022-09-01T11:09:20+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:4d811d67-5565-e442-abe6-e9210aad6c2e" xmpMM:DocumentID="adobe:docid:photoshop:479a7f89-8064-4240-a237-e2c7889a6ce7" xmpMM:OriginalDocumentID="xmp.did:1caa456f-0252-6346-a2ea-2139492196a7"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:1caa456f-0252-6346-a2ea-2139492196a7" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:4d811d67-5565-e442-abe6-e9210aad6c2e" stEvt:when="2022-09-01T11:09:20+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�+y  �IDATxڭ�KLQ��;3m������ą&D�L@W&.4��11>0jԽ	F��Є�t����%qE��
�*}@g:;5-3�C���=������y�3>}�PKHd"+Ǜ��>���ᆃ��/��A(*��tR)+`�>���� -�H. Ĭ�Z0BTuU�� F���F�)�T�6��]�ZUi�i9�H6��=��@V��|�Ѧ �ys�?�:��1o3MP�y�_�`=�6�K��80�{�퀫픩����_=Gp|đ��"�)=]��g
��̋��M��cur�������8�8\ҁ>��f�/��Cc�'���$�$�@��=�/�"R F"�k:(�h�e/��PWCa.�`��pν������[8�q�����^��Z����	�#����j6��iA�l��iz�r:�cj�;�2����¯`�O��� +r��gw�<< w�x$�"��B_�D�K�߸�o�x*D���
X�x)%w�Nnҁ����8��Z�Άx�%e��P<�ݭ]K���X?E/zA���5.�G�|��3���׺h�~��s0:��%l��/��,*�qd!v�_�$�\���T��+����T*����F�Ic��&k�� �^��}���Xq=D�qqAO�b��ݲ+�U    IEND�B`�  Left� Top�   TPngImageListImageList192Height Width 	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:37+01:00" xmp:MetadataDate="2022-09-01T10:57:37+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8ac33e32-9f3e-5048-9d4c-3532138eb0f4" xmpMM:DocumentID="adobe:docid:photoshop:e1d2034c-6c54-f14f-926e-04f6d15de903" xmpMM:OriginalDocumentID="xmp.did:5fa8f5a2-8a46-b542-9d43-49f9de86586a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5fa8f5a2-8a46-b542-9d43-49f9de86586a" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8ac33e32-9f3e-5048-9d4c-3532138eb0f4" stEvt:when="2022-09-01T10:57:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Ǩ�  �IDATx���jA�g�-��̖�^h���(� �E(���g��@|�Ȃ�%PD��荨���Z<������ݙ�͞"���$���������0?h����;7K3#����-����~��ژ��ޚX��s����o��B�Y�^��p�(��t��$�)���#�e������)��un���DL]F�>�3ꦓ��h�/�~����S�)U�*�-� ��Xb�H8�c�~��5����&��@)!kb�᎛Nφ�n��ր��1{�"�+	e��H�v�HO,�%(*��*4���77<���X	k"����)g�Q ��Z@I,��*�� %ԢȜ�wW���$��rq��+��&%dT��3�P�_�B�4)<���`a:2��"Й�E�d.Ml��7�hx�;(�����t�˰Kxgw0jQ��^��p{�h3����M�V���ӊ9!�J�\�w����� �w0$�z��(	\�IP$Lw(R�wL>��_���ܣ�>��`��m[TF�/pg�i=�f�ޔ(�Yph��}D�������`�2[y���L?ۏ>�x�.
��.�!����+{�C�;t�4����ƫ�|�/���rxS��'���@ej��[�\�,8��7��l��<�ߗ��0�;1k�v_���������}3W��a�#�M�X��E��    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
   �PNG

   IHDR           szz�   	pHYs  �  ��o�d   1IDATx���1  �0�_4� ��@�:.      ���xX	     �0��!Hz �    IEND�B`� 
BackgroundclWindowNameOnce Finished - Stay IdlePngImage.Data
A  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:24+01:00" xmp:MetadataDate="2022-09-01T11:07:24+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ceac552f-2eb3-5b47-b3c1-c5ec455c0f53" xmpMM:DocumentID="adobe:docid:photoshop:24a80125-9fd6-744c-8183-cedc9f98d5b0" xmpMM:OriginalDocumentID="xmp.did:cecd1b2a-3619-aa41-bd17-316585b009c3"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:cecd1b2a-3619-aa41-bd17-316585b009c3" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ceac552f-2eb3-5b47-b3c1-c5ec455c0f53" stEvt:when="2022-09-01T11:07:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  IDATxڭW{lSU��sn�mo�u[�uc���HLǈK�H�$>�Fg �D�F>�&J��Є �݀)�
��$&�A���A�l��}Ͻm/m�v���ڞ��s��������"�Զûjj�B�"�T��@!����7���{{.����,J�W� �Y���ǘ�5�pf�0a�aT���*H!�J>٧�TQ�����a�ryN\-T�sf\*VF خًj�z�j�3:.G(��"����)�hr�ϊ@u���cb� ��9�n����OQ"^)@zO�����h;G�?g-���"�l�A�^.�T-�0�m3���y�B�K�P=���80W�L�*�D@Q$���{yt�t��	T�=���}h���ق7�Yᓺ2}�7�¡A����!�ۮ4�}����j�o�V���.���D���~d�o��c��qi���˙)EQ��3�q���e{�]�����Xl}�58=�7愽KQ������i	�Z;[-a��nBـ��<h�<�ʨm��t$͑�~���麦�jZ;{le���QVj��.�e��HP�������9�1�b|ʽ }����Ϸ�"m'3��a�]�y�";.y��ޑ)sT��S�6�s���I�.+����!Mx���X�=|�d���O�'#�2F �B� �5�|7V�C����1`Φ�ko/����a,���85H	�2Ҳ�h���]Ą��U_	����Xj�}�:�;!T�Mp��>Qx��0���Ӑ��	,�Ӏ�	�Ţ��w��Ж��F���!�_+�8#>s�CC�Ÿ�{F��C�13�e�Q�4�`�J@�p����bI���FCa��"�~U�%"=Ѷ��e��ӹ��6�`����ηyI�a0Z�B}�]��g��Y(���r?XK��{�Mc���<��� H���[�O��N(��DBLpN�$�M�C'z����|p#����N3���#> _P��Vow�^���΄w�E�W��V�s�rG���x[��U85���g��y	Dm���D�dB���0�� ����Q�q7t�\�sLU&+!�5��R���P#�����c�	�捿Eu��MN�0>�7�"���z�UB�<V~i���Qp2�.,���{篃/�@]��(�2|J4���~ȃ!x�Z|�d#��L�4��:���EC@,كk/9�ka(uM��㘃R���"�R�Lu�
(Z���/5�>��c��E�W�5�1�yq,&&bc1Ҫm��p5����� ���O�H"	moZ��s&O�4"Jf��[�{�Z�h�s��ڇ`�/�̴�ٝ��ZF�Y��O��u��a���	�ڕw7���+��ش�	D��\@��fM ��v�T�gQ ɷ���QD��Ɍhɜ��Q�"p9�J�)�f��K~�kdR��K+�K[�3�N̡ÖE4R�Ғc��Q��o��@W��<vR�3�ݷ�^�a��Ru1�P�,��H�.�hE	R##$�j�K�$�K���#ٙ��`��=A��
�.03�J�q�ߓ� �t�Lm�%D�    IEND�B`� 
BackgroundclWindowNameOnce Finished - DisconnectPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:27+01:00" xmp:MetadataDate="2022-09-01T11:07:27+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:33024414-1819-174e-baa1-c92e9cddf0ac" xmpMM:DocumentID="adobe:docid:photoshop:59cf1734-3a5f-f544-8e97-0affb646c24e" xmpMM:OriginalDocumentID="xmp.did:03f20825-5636-184e-94f9-484e6711d168"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:03f20825-5636-184e-94f9-484e6711d168" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:33024414-1819-174e-baa1-c92e9cddf0ac" stEvt:when="2022-09-01T11:07:27+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  _IDATxڭ�klU�ϼgv��v��ݲ�B [Kl�,DQ1Fc�"h	��`�� &���Ũ�Q-B�KP	����Rl#�ny����nwg�y�w�;��}P��vv������s�
�;6������ì�((C&JI@Q��{ �;2����+�`�
�������J}������d.��f�=��#0u�����2ud���t�j�װy�>- �����O�"��H� ��"��9"'���u]E����f�*n)/j�#����Kw�	1�e�����2�_� =ڴ��̔ ��)��w�HI������k�GM��p�d"A��p��_�#����9D���a�CG"bZXo^�?�', ߎ�/s�՝'9�*^���������p��ߊ�܇14sõ��/� �6{���|�{2�*���|�)�Vg���Z�{83@��z�W/e���T����=pMu����`��cw���M8���Q�5���������%��Rts�T�s<(�	<��Ѷ�Y�2�MAHk�M���V�5�r~�����ϋr`��iu"���:���g�4Xf|�hV����)%Sd$���O���N�\�o�]��1qF�J,/JN����N�&)�S4&�c�k©���&�M4�Ԑ�7�y$`���}1/.�rR����Y���U��x�^8s�vE�71�� ��L��p�=�|���?��z�b;���D��5ކ�[fף��Y ��+kg��E�P�"ٍ~��6��g��,N�/B�wO����2sWpu�s	|��=�
�^W���w�����<�����W��!P[.u�7����}O����P��C�inp� �l�0°:�g>������C��!�:�E7C�0h����C�b�e'�������@i��·m�nC����}����㕐�gI���-��5o"V�ւ�u����1�w��N>2y�?�o;>~���:��Xm�׼%����sAӍ��?�	(1�ׂ��pDr�\�G����D�c�j���'q>��0�s~��AUi>dB�~x��ŞsFנ����j ��f.�̃��>j��40�������R��k��QO��ʓ��x'T/��������9��z��B�1�p��B��
X�� �"4݊BD6Nu�z!�X���wK-7�dY�,����1�q��88�a$(L#�N�i�]�����e
p��_�F�Ӥ_Qdٹ�R�Z\�ʂ��"A�'h�8'�jBq�p�f4���ri���fe���[�����c�=�+�����}��1��S�5y�T8���I��b��6�]�KhrQ`��N+o���rT1F�'�A�hf�A�P~�Uԏ������j��X�0��2�%����G���L�HO�۝�5�sE1GA�5��ũ�/ut�XY&ym(�]���<Je��]V՘���ި4��8�����Y�`�(�k3m�_K��K-�&��= �����m��D��8:�q������c���Dx
�$j�	����X�#!8�Z��S�ZuW<@ p�^ۮ������}8����?M�w�1B2]    IEND�B`� 
BackgroundclWindowNameOnce Finished - Shut DownPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:33+01:00" xmp:MetadataDate="2022-09-01T11:07:33+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c80d4a19-5922-5343-a254-5f349f3f730b" xmpMM:DocumentID="adobe:docid:photoshop:bed877d9-de31-ea45-9762-b9a2628d2e77" xmpMM:OriginalDocumentID="xmp.did:088575ad-15de-c749-b7da-9019bf33bff0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:088575ad-15de-c749-b7da-9019bf33bff0" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c80d4a19-5922-5343-a254-5f349f3f730b" stEvt:when="2022-09-01T11:07:33+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>Pe�  �IDATxڭWPT��νw�]v�ׂ�yY2h��HkѴ��h+#Q'�����h;��I�T�jM���ZM("�&؆�`e��M4��$T����e�ݽ���{�h"��{�<�������9K0]�sVLJ��5��zB�EU�@2ľw��RU}������m/f���˅��Ч9B^�E��L���'��8*S��
ߘJ}.٥�TQ������ױ'[�' ��8��r��E["$+ 5{Q�_�ڃ���~��S�=�[��[f 1�j1��,��*��sn��?�KQ�C��Ї6e\�����^����3u�?]S56\ �n� {�4/�y�l"�0	0���L�*cbDQ|n���f���ӄ ����� ��`G�e�γB��]F�nhWu;Jۇt6F���1/��� �T���o	����\���%	���1�/\o��Xf�3������.EIbA������t����	v�ئ+���~���3�c)��m��xgJ I��0i�9�Df�<�"�d�\��_Fe.���z���R��+lx2#oJ Ʌ�:[�%IɌ�~4=Kì��Q�"�R�����h۠�qCz����><7 �h�ܥ�ea6I�1��O7�\�{��e�V)��҃�P��IV��t.����~�5��[s��J'Տ�%� �2����<���S�P԰r���V�t��۳Iaؚf�|�W{G&u�2в�s�4`�2'�&Έ���x�g��	e��ҧ�`'!fJX��
oge��<��*�8�FZ�X����0۔@w�iv\|�J~w�,�B���M0��xz���1?�с�X�Y�ވ&�
&�Q�}�x��݈�C$�5�f� p�������}�nU��g,oE5� 	���$��)�&(�d����0
�֮�b�-��t�Ou=Hn�ĳg�C\�9�H,σt6��d}��^����p��#�[��ޞ1�,+����e�D%�D��y��q�E2�O.��Dӄ�XE=Bz[��\�D�]���-���L���=���Ϡ��2tv��Գ(�j�g�i�6����-j�ޢD'�7?�6}؄�=#�ub#)M�Y�(B����[}	���V��0%e�������{��J��A_�ҏ���4�*�LV���~�GK&�/�G�8�2���Z��T��~�iQ?��ن�Cpг ����g�/�鎃����	:2���h�is+��s�} �> ���V��N�_"��F���j�N��
�b���@�ww���x���ۿa<)b�:t�-�"Ƴ�b΋�0gdc����������y#��L6�b2�<���=8��vb^�0w>z������ �l��s�>��� �%�5�M۾��o�Jg�/p�MV�Jx2i���%HM�":�D��cs2��acN\q�n��Ì �mr5�����D,Z:=ީo���-�޼LƉ���1�n���{�A|��9� "����c#ݎ7{tS�k�F �(ns��[�h��y���~ �8>���"��3��С��WZ��}|��K��{�jx>����Qҫ�h�f�ʜ�Qγ-�F��1��O`�V�H,��s����l�臥�ٿ� ��`u������G1P�k4}��բY(�MBI�D[�ѫl��?�S�J��s�z&�mH�E�c�`��~���ihi�p�uͬ�Y�>���2�V�ra;��}#���[G�/DbJ&��>˗V���6���,�ח^�f���H�!UF��6�#���`�&�K=��~uz�)B��+�f���@����P�`��႘,KVA�J��}�up���9���6:8
7��e�r�6~� �va�EI|��dᬒ����OfǶ���n��7e�]~�S3���`�]�V��̀�P)��4!=,.ʊzj�S>��k�7�����    IEND�B`� 
BackgroundclWindowNameOnce Finished - SuspendPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:30+01:00" xmp:MetadataDate="2022-09-01T11:07:30+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b9d4348b-7b47-dd4c-81c9-7317fc2d424c" xmpMM:DocumentID="adobe:docid:photoshop:b6d93b88-5e18-3c4e-87a3-915de2f830ce" xmpMM:OriginalDocumentID="xmp.did:59d422ff-c49e-a44b-80f3-621268e98694"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:59d422ff-c49e-a44b-80f3-621268e98694" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b9d4348b-7b47-dd4c-81c9-7317fc2d424c" stEvt:when="2022-09-01T11:07:30+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>@��  kIDATxڭWPTU��s�݅U �E{�##�S��cjN��#�Sj6�6�3���TVf��9��gi�Z����$�R1Y`w��� 层�{��ι�n�`?��=������������-�)C!�9YD%1 ���� $����v[�a,�B;�k��Q1�{ǩ<�}*�</GH�^�x���9�@UT�T�v*NU!��V�ŢA�#�l�3��+��8C��H������]v����+.��*�=�[��H0�<;�z� $m��ɉ�C�Π�(
>���������j���C�8r�ϴ	 ;9'ȅ�.aᲁG[�C�NWTƆ�x�5Lp��'����Kj��c$z�Ǖ:�C�2Q���������	@��3�0�Ks|���γ:�*�������w�Vc�~��V�e����ZJ��	sk�Թ?g%��N�6��:_p�v�f����Rkl�咶^&�) S[c��%�#��圹�����kk�4E�W�釂�l/���7K\[�w5�؝�2����N�-(o���H�R���@������"�\�Ծ"�F�M�{F����Ai���A�Ĵ���v���-,�c'i��g�LX��ٿ���
l��	X�Ҍ`�Ҟ���b���ҹ���Ǆ��
�ASo��(*iQ?.�
��@D<c ~��4���w����M׫@+��}̴DazR��)g�������R�0;�-���O��wRM:m�^�Z�n�>	���������/�7��"��O��Y��Jm1�]�um���f=�b�:��u&џkҺ"�C��
�K7�����^��3ᝠ»�z���+A������a�ۯ�$n).��]�X��Ga,�歷x�av��>z7��Z�6��~���uNm|܈�0vē��3�	�q�.��v`��8�5�)����*+-�� �*�!Fo	K��ܧ9�1�x�w�-(_��;gf�cɻ�18��lM��s>��ϔi T�Շ1�}l+xC�����d�O�죓,bs���}�s�
�V�CY���0 �$�X��K藑�<�����X��4�Vl�ZR"��p)Q2
��@�*?N'aSf��8H��ιr*8J��A�m��tl�T�����0h�:��A�f� �
uh�Ū2T�5 ����3n�W_���e�*���!E7sr?̞�t��7�bK>cdu`G$�G$�`��@�0�6l�,�vyH =��j����K+0z��YQ�=!/��"�$�h���"�,�H�\CH z*��
�W�B���l���]qr�4�E�9�r"	&�s��`X�Sߟ �Cw�:Y@������v���L����^�(Y!�BC���5b���B`�W`��-���� BXrJ�F�r�j��21wڀ��U�N�u�X<׷@R��a��5�}���^Ct�1���4�T�ã��v`�=%�*�~�s������}������VF�����#�X,=xQ:�Յט����Cz5��Ш`����"0���/-��׀D������K�>iL:r^�@�����Jy5r�l���9TܭcS�P�؋�s5� �n))�$�[
G3#��(d��a���� >����d,mB����XNB_�KJ�?���ݽ)�"    IEND�B`� 
BackgroundclWindowNameSpeed LimitPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:46+01:00" xmp:ModifyDate="2022-09-01T11:07:36+01:00" xmp:MetadataDate="2022-09-01T11:07:36+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:564817a0-ba0b-ff46-8e0d-3e3684c4a162" xmpMM:DocumentID="adobe:docid:photoshop:6755485c-4eeb-e341-90d6-19acdc5d0ff0" xmpMM:OriginalDocumentID="xmp.did:b6a41e6d-297c-0c41-bb28-86cc694cb847"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:b6a41e6d-297c-0c41-bb28-86cc694cb847" stEvt:when="2022-06-27T15:59:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:564817a0-ba0b-ff46-8e0d-3e3684c4a162" stEvt:when="2022-09-01T11:07:36+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>2W�)  �IDATxڵWPT����DyYlb�4�)��P\e��J5FL�v�щ("/E��F35hhj��4
8�F@�UPc�
b������}��H���ٻ������;�O�9Whh��L�2J�̲��WTT�?�9�p��̗Qѯ�Kh�
�9DA��B� ��3������� [6��3D�
�Ba�嬙���.�~�9r�����<lj���7�����Mf�� �L�p)���=/ Z�<���4ovͪ8��ys!�Ɇ�@��pX��?.�t���'OZe���*-)��� ̚�\�5�>M3t�[o��^���d�׷��M�w+�>n ��
�@�=�xO�bR�CA����9��P̟�$_�9�B���uu�=?
@T�=��P*U3�S�����	���r�<���a�$ `��w���h�z�h\�q{���M&S}k�D ��*�Zw(������*�S����P�P����N�C����9P�X"���m�f��XXZR�bH aK#��dLf֞]L�����0V����ەڼ���d(���[H߽�cY.��ˢ? ��F�ug��5tlLm��ݕ;��u:�vy@,� Pnc@Ԁ�h&�qƚ�`5����5�d��p���?s��,���Ң�N G��2��'����)S;�ű(�t�hh�	CC� fJ4��"�E��d�$y�+��"��d zB��{�W�]=�a�Ó�֒���� ��"��
�)1�]j���`�`�_Dp��5Mj,���o���E*7Q�U��'�~S��#����G9{ԫ����j�X�͂_yy�#	��p��R��YA�Bfn��,�W1����[�R���_���h���Z' v����Gϧ;��@<#g�gՂ፵�0'���0W��Еϝ<g�����y�7r%��.��/:���446J�D2Z�`>bb�@�� �^0�F�;ܣ{V/�	�F�!o⽼C�W�^�.-)�X����u��Z-�k[����P�6/DC�Յ��4<|��[B������Uq���'/��Ty��t[2
`&σK§(�{%>>u���b���j= S�gf�c�ԩ����y(%�@�w��OR���F@�����y�4~<��f ��܅>9D:G@�לZܾ}���H�=�����2J�x(7���A�,k��/*O)��wSv&��`08�(8�IoU�Ca�Ƴ� �0�8݌��f�HJ& �	 s`��?d��"2����heol�{CC#v��$+��2e2R����`�F����y$Hڙb`AFz*	A �7׃24[�J��#��~N�ec�=T]��F�(�n���-G������?R��p=|�����ﷆ����Ŀ�8,���;��n�y�:��# `��z=e��!'�g1���Y���K�η&����~5g����_B�r�f
��E�����_�NBI\޵y����U�̈́\��?8�]__�[�")	�<�B��}�H�a����[�Z�YZJ�өd�!�@�W�цM�Yz��Nś7m�����n=ų
��w�^8���jg�>�i��;��qݿh%d�3q��;��3�/#o/ψ����#l��ATb����S7����W~��V2Sh ˨$����dC[�S�˨�u��L��%�\��a����K7�� 4l=��8�p?�uG@MAYY9���yR~S\�}���� Rی�XՋ?j�^�i��H�H^n�r���mI-�u{v�+||F���y�w=~�{3�H�I-��2à �4��W6mܨYn�������f�yxM���-_�Z,M�0�LCò־xr�VVV	�Ν#�����X�H�.///sLT�f欙`Hk�z�q���q�BaO[[��@I#�Iv_�����f
��2m�tˤ�]ƌ�\ݬ�a�^����h�{���͛r���fN�i8��p�~�)�p*��ӡ�8�C��R��������v:2\(    IEND�B`� 
BackgroundclWindowNameDownload in BackgroundPngImage.Data
�	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:57+01:00" xmp:MetadataDate="2022-09-01T11:07:57+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:74cd029f-22fd-4343-a26a-0f034390f58c" xmpMM:DocumentID="adobe:docid:photoshop:85e04310-3a95-f643-8199-5af10c9b1696" xmpMM:OriginalDocumentID="xmp.did:69da3e75-e159-464c-9549-280c60220390"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:69da3e75-e159-464c-9549-280c60220390" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:74cd029f-22fd-4343-a26a-0f034390f58c" stEvt:when="2022-09-01T11:07:57+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  �IDATxڽ�]HQ�߳3�i�XQٯD�ETD���M7]E�V�֍�7^TwIaQ]DB��RA�AY,eijV�Ϧ�3��9�������̤~����8���=�K�Ν����B@)---)>g��? �{v��w��UȲ�p8l	1) ۷nA]�CK�I}ݿz,!&@�ĸ ��Vk"���%c�M�$I(ܲ�fΰ/�(�`��4�t]�g_�c� �����
6��Ą �I�/B�	u 6�c9�
�M�cI�I ��X�^w<D����*���;/�&*�f��~��5�rC�s�J/BEI�s �I����4�g� <i�>L���B�/�Whv�t�ր��z��t 29��o���E"�?a�@�)���Du�h��ڵ�7})N︇t93��ĥ�h�n@��'�F�E�#�=�z���M҇X7�IՐ��H뛉uR���'!c�2*n
�24@i�������W8�� ��D��'��F�0�\�I	��)ĵ�)�tu[���][$��5jZ+�>g$�i��q"��/�F���Lm��ܽ�|r���b/W�}R��5�r����	���W��ͧ�Ƌ'�u�u�-tM}o6�b1i�+�����(��4���G�!�0�b-�ځzZ��C�YYja�����P{Qrs�W�W�8�����(�]W�#�~���:�.�
2���N�P:=!��|Rz�7<��и8�ޗ÷8=���p�@m������3�^�n ;p�i>�w����^�n!�]�`^3�A�F｡��-����R�P�}������ l��j�U�^1f!.2���ѩ
��z�A�������:�E�?�@0����*���#(���ŧ�S���Uk! m#Tkk,W�����v�,�&    IEND�B`� 
BackgroundclWindowNameUpload in BackgroundPngImage.Data
�	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:08+01:00" xmp:MetadataDate="2022-09-01T11:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d785d370-05ac-8c46-9266-34272c48ae57" xmpMM:DocumentID="adobe:docid:photoshop:698042e2-1780-5c40-93fc-52fa2955f328" xmpMM:OriginalDocumentID="xmp.did:e2bf7891-7e9d-8a4d-9337-84fc89c4569d"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e2bf7891-7e9d-8a4d-9337-84fc89c4569d" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d785d370-05ac-8c46-9266-34272c48ae57" stEvt:when="2022-09-01T11:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  �IDATxڽ�oLeǿO{w�hKVa	��${a�!Q��!N^���B���?����{�M���h��7K�e�EEͲ-[�6�����z��]{���T��X�G�4�������>-g���u3�!�4mp�����p��keם��kpUU!v��p/~���bW غ�p�b� �AT���ot���7��� f�n���boy�<�x���Y�<kz&��u�ƪ��>}��z����7�GV�-L쨁¦�3a	�J�u]/Y[��Mg�11�����2nGҸ���7������u�ݦ�AL�Ux�u���v,���Ő�mpB�������� ��6pg2����#3�8un~��苸�\4��˽���m$���]�?�.WP�tY��å&ȍ^�?���;���Z|��X�����D� l
���=�>��U'���cb�j"�&�h��.D��y�i嬈�V�	Z�D2�t�2`d�h���ѽh�i���!nLEqC�_5S����n������� c�o��A%5�ᨊ��f�	5����Z���f�JY�O������6���K8�������%Ǎ=m�vHa+�k�&�{��mxg���6����Õ�V��ʾ���V��!�%�/�!�t�[6������;X��i'P�o��lL���&����y�ȵ����G;?�d ��u��͕hg�+��YU{E�:����If��p#��zU횬� {r^�;^��9�`����)���RzSiWƺ����W����3,�r�4�B�譩t҅O��������O <Z��y�iOe��.f3[�@��q"�A���R	�!24��|������x$'>[��>7����������n���j�~�J8� .vvV��jz    IEND�B`� 
BackgroundclWindowNameSkipPngImage.Data
:	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:14+01:00" xmp:MetadataDate="2022-09-01T11:09:14+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:32cf113e-1248-bc44-a71f-672f26c5d91a" xmpMM:DocumentID="adobe:docid:photoshop:57ffb0f6-9680-5349-ad59-8e90e59ef86a" xmpMM:OriginalDocumentID="xmp.did:b19fb083-9f64-7747-84c2-653ae1e8dccf"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:b19fb083-9f64-7747-84c2-653ae1e8dccf" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:32cf113e-1248-bc44-a71f-672f26c5d91a" stEvt:when="2022-09-01T11:09:14+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>1�bm  IDATx�͖KLQ��i)h�B	hh	PP7*1�-�@D6|`A )ĵ4qa"�	[QP_]�BA|�ZTwP4.1��$l{�eh;3tڹP�'i&'��w�s;)G��,���u+$��¶��a�E4[��P����^������v��@D������ �
@��:]LQ���n���! Ķ`����0�nmi�l��Hv| ܶ���e a}^x���i�5�CȽ�O"����g_������#�dZ���	�L5�W�2P7&8@X��6tk���S�xWN����d�v��� GpQ�����jr�WA��_��ڑ  �X����8B�|]��$k�#`H�H�����,�	��,�u��������1��~P�@0}���I�G}n'2��� (Rl��)�5xj�_"���L�����/�������%����X=.�	{�3 p���a�RIv8ҭ� �p��H]>�Y��[������]S������=/!ן�.^�y�%����1IH�dN���s��r���Լxt\��wŧ�Sǣ��SF3����@�k	@�BN��n놠P=���+R��}� �������1�=i	{�z������
�Z�+���JF�� �����oFuN��zi� �$ �, �ىyh��	c�!ȕ��K�H �M��vL��*��q�$���?R �h� �J�:=�5�8�� ��7q����LGL�Ԗ 8���l�KOY��uf`}$�[�,�!�D    IEND�B`� 
BackgroundclWindowNameDelete in BackgroundPngImage.Data
w	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T16:00:54+01:00" xmp:ModifyDate="2022-09-01T11:09:21+01:00" xmp:MetadataDate="2022-09-01T11:09:21+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:1758d269-8c01-104f-a653-e35e4ea393dc" xmpMM:DocumentID="adobe:docid:photoshop:1b5fbac2-806b-ae4c-a4fa-5db1c57fb8a9" xmpMM:OriginalDocumentID="xmp.did:ecd867b8-9017-d948-b067-f3c9ddfbbd1d"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ecd867b8-9017-d948-b067-f3c9ddfbbd1d" stEvt:when="2022-06-27T16:00:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:1758d269-8c01-104f-a653-e35e4ea393dc" stEvt:when="2022-09-01T11:09:21+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>� s�  TIDATxڽ�KLQ���1���R
�B4h�6��*�J����&&&�5Q�B�ƅ��]��+	+�mL(�A�Z�����w�g��3C���&�������gZr�����7�޻t���uA ������}��!Y$��i ��albR�i R_l9���T ��!� ������w�ɁeЛt�{�().�/A��k��h����Ku,� R�'���~�ΌN ��S�NԁԤgr"'�l��a�<�(dҵ�S *�����m���@�IϻjIg��B���?{�ɼ������x���(�M�����O�B�� ��p:��H�헁�Dq���-��T�nԪ��y �P���3L{����);������ԉ���ėb]��E��g����A��I�������pIt�E��nw���8�!�!�ِ���A���q/ج8�"��NX���m�Y�4�jw��3Ӌ!V�:��h:��-~��تpϱ�������c��\5u[�``	Q�*.�"�)�r y�J�Z��k�BQ������c
qU�\P&]��@U�A^��E�
�9���k�
@d�o/�: rq@J�t-�� �	���F��s4�֓�4�P@�Ł�Q��1��
��.0����z��R!�������q\*7��_b�!�GkOu�v@�qwO��fpU���E1,�yˤ;j=���>�on�rXb�h6�Ӭ"lD5a�&�WE	����9�C��n���H����������IM<�l�N��$ �&��*��ޣD�	��4Ӫ%�
a%�N��_���]R�j�����    IEND�B`�  Left Top�   TApplicationEventsApplicationEventsLeft� Top�    TPF0TPropertiesDialogPropertiesDialogLeft�Top� HelpType	htKeywordHelpKeywordui_propertiesBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption
PropertiesClientHeight�ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize�� 
TextHeight TButtonOkButtonLeft� Top�WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top�WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TPageControlPageControlLeft Top Width�Height�
ActivePageCommonSheetAnchorsakLeftakTopakRightakBottom TabOrder OnChangePageControlChange 	TTabSheetCommonSheetCaption   Allmänt
DesignSize�c  TBevelBevel1LeftTop,WidthzHeight	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelLabel1LeftTop7Width1HeightCaptionPlats:ShowAccelChar  TLabelLabel2LeftTopNWidthHeightCaptionStorlek:ShowAccelChar  TLabelLinksToLabelLabelLeftTopeWidth,HeightCaption   Länkar till:ShowAccelChar  TBevelBevel2LeftTop|WidthzHeight	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabelRightsLabelLeftTop� WidthBHeightCaption   Filrättigheter:FocusControlRightsFrame  TBevelGroupOwnerRightsBevelLeftTop� WidthzHeight	AnchorsakLeftakTopakRight Shape	bsTopLine  TLabel
GroupLabelLeftTop� Width$HeightCaptionGrupp:FocusControlGroupComboBox  TLabel
OwnerLabelLeftTop� Width&HeightCaption   Ägare:FocusControlOwnerComboBox  TImageFileIconImageLeftTopWidth Height AutoSize	  TBevelRecursiveBevelLeftTopBWidthzHeight	AnchorsakLeftakTopakRight Shape	bsTopLine  TEditLocationLabelLeftZTop7Width%HeightTabStopAnchorsakLeftakTopakRight AutoSizeBorderStylebsNoneTabOrderTextLocationLabel  TEdit	FileLabelLeftZTopWidth%HeightTabStopAnchorsakLeftakTopakRight AutoSizeBorderStylebsNoneTabOrderText	FileLabel  TEdit	SizeLabelLeftZTopNWidth� HeightTabStopAnchorsakLeftakTopakRight AutoSizeBorderStylebsNoneTabOrder	Text	SizeLabel  TEditLinksToLabelLeftZTopeWidth%HeightTabStopAnchorsakLeftakTopakRight AutoSizeBorderStylebsNoneTabOrder
TextLinksToLabel  TEdit	GroupViewLeftZTop� Width%HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNone	MaxLength2TabOrderText	GroupView  TEdit	OwnerViewLeftZTop� Width%HeightTabStopAnchorsakLeftakTopakRight BorderStylebsNone	MaxLength2TabOrderText	OwnerView  �TRightsFrameRightsFrameLeftYTop� WidthHeight� TabOrder  	TComboBoxGroupComboBoxLeftZTop� Width� HeightDropDownCount	MaxLength2TabOrderTextGroupComboBoxOnChangeControlChangeOnExitGroupComboBoxExit  	TComboBoxOwnerComboBoxLeftZTop� Width� HeightDropDownCount	MaxLength2TabOrderTextOwnerComboBoxOnChangeControlChangeOnExitOwnerComboBoxExit  	TCheckBoxRecursiveCheck2LeftTopLWidthwHeightAnchorsakLeftakTopakRight Caption/   Ange ägare, grupp och behörigheter &rekursivtTabOrderOnClickControlChange  TButtonCalculateSizeButtonLeft/TopHWidthPHeightAnchorsakTopakRight Caption	   B&eräknaTabOrder OnClickCalculateSizeButtonClick   	TTabSheetChecksumSheetCaptionKontrollsumma
ImageIndex
DesignSize�c  TLabelLabel6LeftTopWidth9HeightCaption
&Algoritm:FocusControlChecksumAlgEdit  	TListViewChecksumViewLeftTop"WidthzHeight;AnchorsakLeftakTopakRightakBottom ColumnsCaptionFilWidthd CaptionKontrollsummaWidthd  ColumnClickDoubleBuffered	MultiSelect	ReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder	ViewStylevsReportOnContextPopupListViewContextPopup  	TComboBoxChecksumAlgEditLeftZTopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeChecksumAlgEditChangeOnEnterControlChangeOnExitControlChangeItems.StringsXmd5   TButtonChecksumButtonLeft� TopWidth� HeightAnchorsakTopakRight Caption   B&eräkna kontrollsummaTabOrderOnClickChecksumButtonClick  	TGroupBoxChecksumGroupLeftTop"WidthzHeight3AnchorsakLeftakRightakBottom CaptionKontrollsummaTabOrder
DesignSizez3  TLabelChecksumUnknownLabelLeft
TopWidth� HeightCaptionChecksumUnknownLabelShowAccelChar  TEditChecksumEditLeft	TopWidthfHeightTabStopAnchorsakLeftakTopakRight BorderStylebsNoneColor	clBtnFaceReadOnly	TabOrder TextChecksumEdit    	TTabSheet	TagsSheetCaptionTaggar
ImageIndex
DesignSize�c  	TListViewTagsViewLeftTopWidth~Height� AnchorsakLeftakTopakRightakBottom ColumnsCaptionNyckelWidthd Caption   VärdeWidthd  ColumnClickDoubleBuffered	HideSelectionReadOnly		RowSelect	ParentDoubleBuffered	PopupMenuListViewMenuTabOrder 	ViewStylevsReportOnContextPopupListViewContextPopup
OnDblClickTagsViewDblClick	OnKeyDownTagsViewKeyDownOnSelectItemTagsViewSelectItem  TButtonAddTagButtonLeft� Top� WidthPHeightAnchorsakRightakBottom Caption   &Lägg till...TabOrderOnClickAddTagButtonClick  TButtonRemoveTagButtonLeft1Top� WidthPHeightAnchorsakRightakBottom Caption&Ta bortTabOrderOnClickRemoveTagButtonClick  TButtonEditTagButtonLeft� Top� WidthPHeightAnchorsakRightakBottom Caption&Redigera...TabOrderOnClickEditTagButtonClick    TButton
HelpButtonLeft6Top�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  
TPopupMenuListViewMenuLeftTop� 	TMenuItemCopyCaption&KopieraOnClick	CopyClick    TPF0TRemoteTransferDialogRemoteTransferDialogLeft(Top� HelpType	htKeywordHelpKeywordui_duplicateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionRemoteTransferDialogClientHeight� ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize��  
TextHeight 	TGroupBoxGroupLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize��   TLabelSessionLabelLeft/Top	WidthMHeightCaption   Mål&session:FocusControlSessionCombo  TLabelLabel3Left/Top;WidthhHeightCaption   Målfjärr&sökväg:FocusControlDirectoryEdit  TImageImageLeft	TopWidth Height AutoSize	  	TComboBoxSessionComboLeft/TopWidth�HeightStylecsDropDownListAnchorsakLeftakTopakRight DropDownCount	MaxLength� TabOrder OnChangeSessionComboChange  THistoryComboBoxDirectoryEditLeft/TopMWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxNotDirectCopyCheckLeft1TopjWidth�HeightAnchorsakLeftakTopakRight Caption#   Dubblera via lokal &temporär kopiaTabOrderOnClickNotDirectCopyCheckClick   TButtonOkButtonLeft� Top� WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft"Top� WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftxTop� WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TPF0TRightsFrameRightsFrameLeft Top WidthHeight� Font.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 
ParentFontTabOrder OnContextPopupFrameContextPopup TSpeedButtonOthersButtonTagLeftTop2Width+HeightCaptionA&ndraFlat	OnClickRightsButtonsClick  TSpeedButtonGroupButtonTagLeftTopWidth'HeightCaption&GruppFlat	OnClickRightsButtonsClick  TSpeedButtonOwnerButtonTagLeftTopWidth(HeightCaption   &ÄgareFlat	OnClickRightsButtonsClick  TLabel
OctalLabelLeftTopNWidthHeightCaptionO&ktal:FocusControl	OctalEdit  TGrayedCheckBoxOwnerReadCheckTag LeftATopWidth"HeightHint   LäsCaptionRParentShowHintShowHint	TabOrder OnClickControlChange  TGrayedCheckBoxOwnerWriteCheckTag� LeftgTopWidth"HeightHintSkrivCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOwnerExecuteCheckTag@Left� TopWidthHeightHint   Kör/ÖppnaCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupReadCheckTag LeftATopWidth"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupWriteCheckTagLeftgTopWidth!HeightCaptionWParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxGroupExecuteCheckTagLeft� TopWidthHeightCaptionXParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersReadCheckTagLeftATop4Width"HeightCaptionRParentShowHintShowHint	TabOrderOnClickControlChange  TGrayedCheckBoxOthersWriteCheckTagLeftgTop4Width!HeightCaptionWParentShowHintShowHint	TabOrder	OnClickControlChange  TGrayedCheckBoxOthersExecuteCheckTagLeft� Top4WidthHeightCaptionXParentShowHintShowHint	TabOrder
OnClickControlChange  	TCheckBoxDirectoriesXCheckLeft
TopfWidth� HeightCaptionAddera &X till katalogerTabOrderOnClickControlChange  TEdit	OctalEditLeftATopKWidthFHeight	MaxLengthTabOrderText	OctalEditOnChangeOctalEditChangeOnExitOctalEditExit  TGrayedCheckBoxSetUidCheckTag Left� TopWidthMHeightCaption	   Sätt UIDTabOrderOnClickControlChange  TGrayedCheckBoxSetGIDCheckTag Left� TopWidthMHeightCaption	   Sätt GIDTabOrderOnClickControlChange  TGrayedCheckBoxStickyBitCheckTag Left� Top4WidthMHeightCaption
Sticky bitTabOrderOnClickControlChange  TButtonCloseButtonLeft� TopbWidthPHeightCaption   StängTabOrderVisibleOnClickCloseButtonClick  
TPopupMenuRightsPopupImagesRightsImagesOnPopupRightsPopupPopupLeft� Top; 	TMenuItem	Norights1ActionNoRightsAction  	TMenuItemDefaultrights1ActionDefaultRightsAction  	TMenuItem
Allrights1ActionAllRightsAction  	TMenuItem
Leaveasis1ActionLeaveRightsAsIsAction  	TMenuItemN1Caption-  	TMenuItemCopyAsText1ActionCopyTextAction  	TMenuItemCopyAsOctal1ActionCopyOctalAction  	TMenuItemPaste1ActionPasteAction   TActionListRightsActionsImagesRightsImages	OnExecuteRightsActionsExecuteOnUpdateRightsActionsUpdateLeft� Top TActionNoRightsActionCaption   I&nga rättigheter
ImageIndex ShortCutN@  TActionDefaultRightsActionCaption   Stan&dardrättigheter
ImageIndexShortCutD@  TActionAllRightsActionCaption   &Alla rättigheter
ImageIndexShortCutA@  TActionLeaveRightsAsIsActionCaption   &Lämna oförändradShortCutL@  TActionCopyTextActionCaption&Kopiera som text
ImageIndexShortCutC@  TActionCopyOctalActionCaptionKopiera som &oktalt
ImageIndexShortCutO@  TActionPasteActionCaptionKl&istra in
ImageIndexShortCutV@   TPngImageListRightsImages	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
	  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:09+01:00" xmp:MetadataDate="2022-09-01T11:02:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5b7adb81-36dd-bc48-ba23-0569e2550d2c" xmpMM:DocumentID="adobe:docid:photoshop:1cea56de-8eb2-034d-aa4f-b5ce08fc08b1" xmpMM:OriginalDocumentID="xmp.did:bd819090-28bf-b349-89cc-8656a2332f78"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:bd819090-28bf-b349-89cc-8656a2332f78" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5b7adb81-36dd-bc48-ba23-0569e2550d2c" stEvt:when="2022-09-01T11:02:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�}��  �IDATx�u�[HQ���n���Z�����c%��E���YiL�03�%5$$J��z�-)�ijiꦮ��`dQ$����e����:�Lg-F���o8s��|�}3��(,��0�l-[(�@		�	�*z'���O���	����u����n$��E�F����������@qq1�!��%Ű�,�6J��e<�$�E�_&���ៀ��5�R�	K�eB�R�w�
�+��2(�D	]��4eI��O���^���{ң�I��/��ç�	`W*��%�U+��lljf�	D!�{������-���=������x�ݽRv�8��2Muaf�5�5R���}g���A�y�Mq����:��>��l�
0�'�J�`.�>|��^_o/�� �od����xx��!J����D�b�=��O���ˣ���]`��?�t�KBD���}R���m�(J:B�?���7�� �#�pNh�=~Ri����sx]Ӯ�`#T�P��9�P?nD,������'�d��3�wT�M�`��������[[p��Ah��iѢ�!���,���Rw'm�V������
�moG����7X���� <��r&wfg%��0WAeu-�@�	B 0��� ����.���L(��
�߿��zGfF=�kT�qE�O}z���� ����LD�!�"R�uPs�B�W_�E3��a���=�������죜b=�vܩ�V\[�ؗ�E6R�$�g�5n��{yӢWL�;���^��    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:12+01:00" xmp:MetadataDate="2022-09-01T11:02:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e9d69505-da96-b640-9af0-aaf7fae84253" xmpMM:DocumentID="adobe:docid:photoshop:fe7bf818-b394-f446-9d05-79810945c22a" xmpMM:OriginalDocumentID="xmp.did:4089a4f6-568f-f14b-9f96-e85fac40ba31"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:4089a4f6-568f-f14b-9f96-e85fac40ba31" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e9d69505-da96-b640-9af0-aaf7fae84253" stEvt:when="2022-09-01T11:02:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>`��  {IDATx�u�MkAǟ�h^v�ڤ���+R[��*i�&h�JA�O`��E�x��Z���֦1/-�ZP���&��m�$�ug�g�twc�������7��0�,�2��H$�
�K	�&�Y��G���o�E��x�ɴ�a�Rz�h�ne���@����h����YD�~<��"��ⲇR҆vmM"]�N���) ���T~�bI"��D��W������B�$%t�$�o
�'3����ѱ�#g��<q��,S��Of�V� x9�L����$�����b����)�*�#>���~ii��c%���g��i��V՘H�����j��m;.�>p����ǕZ�j��p��b�������:��\��V��rwvfU�|vQE��no��4�L�5�Y���l�ܮ�	���
� �`����r9��eA�2�|��z�] K�0��/�/A�T��w���C�B`bـ��� X�&������L2si�~�_�6	z�|^����c8T���H�S����7�%��y5���z `�%�u�WA	!��i�ѧ�5A��XF+�^H783�~�����Z�v
C���P� ���C������U�R�
�������� w    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
	  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:15+01:00" xmp:MetadataDate="2022-09-01T11:02:15+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:759cc3b6-0b75-3642-a75a-d9a08a216678" xmpMM:DocumentID="adobe:docid:photoshop:63b9f3be-b620-be4e-90be-09693bb62be4" xmpMM:OriginalDocumentID="xmp.did:c7d3454f-790a-0c44-8f38-27b9c04bd6a9"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c7d3454f-790a-0c44-8f38-27b9c04bd6a9" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:759cc3b6-0b75-3642-a75a-d9a08a216678" stEvt:when="2022-09-01T11:02:15+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�� �  �IDATx�u�[HTA���͵�U�hwE"�H2(��e��eYJ)%*A=�/�CB��D/Q!	����y�mW�������%�����v�9�gf�]�f��0�|���c�A�p��-�8H		V�,yf*srr~a�����k�4��R�H�DF'y���:��_�f���K��I���<�:	%��5�R��G�W!{�O��^�;_eS��dE!$��Ѵ��o嵵F����#/7'uY๣����,_�QF��3K}��� Z����O�x��?@���'$�\�<z��B����1?$�b�Z�\�h��]6�����7j6o��C#���a��s���,޾�=cD�:�罊�&��i��gzm86�%a[䱔��,�
��wH�,kMfzC ��:�0<m��w �<@,;��a�H�@w�
���K�$k��恒����A�&��*��ہ+[��y��w��� ?B�=� E�=kvʁ���`�nm�^����c�_W~ 3���%"*!�q�hB��<
�o���t��a棆�@]�s���ޑ��i��އ�G�M���Ƶ�L���=�S���Ik���� �2\�>��K�ל�|�Թ?��4>��JT��I�(Ib��c((�W�_
�B~B&����*��3L�~��U��g��D�x
B�(��s���_ &���T����dŽ2Dc`�5;g��)�f�;��5��M    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:18+01:00" xmp:MetadataDate="2022-09-01T11:02:18+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:1a7ecbed-839e-604c-8404-8b59e2d7ac03" xmpMM:DocumentID="adobe:docid:photoshop:4a05ce76-501d-014e-a4db-548903bf8baf" xmpMM:OriginalDocumentID="xmp.did:662c693c-a43f-bc40-8d18-5618731047ce"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:662c693c-a43f-bc40-8d18-5618731047ce" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:1a7ecbed-839e-604c-8404-8b59e2d7ac03" stEvt:when="2022-09-01T11:02:18+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>I�̮   �IDATx�c���?��Y��3`��@A����#8 H/#̀��X�9�3���|���'.C�����}���4 	��JOf%� tÀ0�5@BL�a�y`���W3���i??�lܴ	�!=%��ū7��3X ���b�,�c&+-�#���@(f2ӒX�02b�ô�s	�� F������0M����i��t��A� �  ��o^    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:46+01:00" xmp:MetadataDate="2022-09-01T11:02:46+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8aaab8fd-fc79-4640-b723-6ad8c761b2fa" xmpMM:DocumentID="adobe:docid:photoshop:0bf49fb8-5154-3648-9847-bebd7fedb212" xmpMM:OriginalDocumentID="xmp.did:27ad1779-668d-4044-9331-a61efba7ca17"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:27ad1779-668d-4044-9331-a61efba7ca17" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8aaab8fd-fc79-4640-b723-6ad8c761b2fa" stEvt:when="2022-09-01T11:02:46+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>s�Z   �IDATx�c���?��Y��3`��@A����#8 H/#̀��X�9�3���~����.C�����s�^��4 	��JOf�k�����9���)I>ޞ(�`�k��M�6�_�����6���[���A��0x�����JK:'!1��̴$f�����0m�\�14���b�d@ ć2Y.��D� =@l�\�@ �  �	�:���    IEND�B`� 
BackgroundclWindowNamePaste rightsPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:48+01:00" xmp:MetadataDate="2022-09-01T11:02:48+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8e4e0077-43d7-614f-b817-c5a9c863b158" xmpMM:DocumentID="adobe:docid:photoshop:509e1619-7cf3-4b46-b822-cf94ed6d3915" xmpMM:OriginalDocumentID="xmp.did:f3af905d-f299-1249-a8be-3af395de2041"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:f3af905d-f299-1249-a8be-3af395de2041" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8e4e0077-43d7-614f-b817-c5a9c863b158" stEvt:when="2022-09-01T11:02:48+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��1i  �IDATx�c���?###2��G���?c���l�ϋp �^q�������$��ʫ$(Ȼ����\��+?���|�·k �?��t1|�0�D�O �$h`,��ʯ��R����s�C{3���;��i�v������j`$���-
��������O;�>c�������{�+�:��L���A��eB7�XĀ� �p�A���X8҄i�ٹ� �ӏ����u�P8Ԁi�-��)��(̙�������_�|�����8P�j ����� ?o��;�|���{VZ���}5��W��t�j��?~0�D�2,����̴$f��=U������]4�l��
Lk�� �\7`G�O�Hp���0��	.�R���Q ـ�z$� =;����s�3   W^��J*�    IEND�B`�  Lefth  TPngImageListRightsImages120HeightWidth	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
�	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:10+01:00" xmp:MetadataDate="2022-09-01T11:02:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b987d3a4-576c-0841-8a26-bd069158cda6" xmpMM:DocumentID="adobe:docid:photoshop:ace24ca5-9841-514d-a778-5c201fae19d2" xmpMM:OriginalDocumentID="xmp.did:18550348-d9e3-6245-9980-dcc5f553dc98"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:18550348-d9e3-6245-9980-dcc5f553dc98" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b987d3a4-576c-0841-8a26-bd069158cda6" stEvt:when="2022-09-01T11:02:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  �IDATxڍ�mL[U���RZ��f뚾PNc����q����hXY��7��D?�L?����03��n��/qn�׬c�"]�X	�1~-ݠHCKiｽ��빷t��pO�{�y������s��TUE�8���̼����&Y�|>_�� `ww��+5���4RJ˘��-Br��;w�����P(T�i��~T�*�B��j�y(`o_��P��`H��U�y��˷�s¼������U��ޫ[����Я�}mmmJ�Oǅ��RU�B��~ָo��{B�O���hTE������/�lǅ?Y962CM�n^�����J�LRr�k/�]��g�u�'��b�N5����@���peF�/��*�ɘq��G��؝�~A�r���;����[xc�(Jf��8b�w�P�Q���U��Y�jj�]�ܠ��p�N�S-zVx����غ�y�2`82��2g6[�r9�`T�`�� ���d�= !����wf���{����z�.�K����pk�܍`s���o��݀Db���~���:��<}wn��Y�9=C�ۭ��4�jj���#��0!:�@i:�d*	����׈�Xb&�����������<�Fn�ė���nA���D\�N*=���g���̫/�T����^C�Z�����~|r���-p�[�u��D�sկ�֝��زE��_f�8��z/Cmmo�G,Cm�A�7�Q�.?n�_���u+;:�y�VM�'�ᒭ���=��;������v��'Ŵ���-�|��N�$�z=�@����݇��L�H�nA*5o�*�S��A��墿�tVXK�2M��~6P��G��dښ�J����%��&<Ǖ���I���m�Ͱv6)r��(��M�ʌ�Ȅ��I[WjKK��1��?�R}
UG�    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:12+01:00" xmp:MetadataDate="2022-09-01T11:02:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:03d57e26-91b7-5440-a88f-df46974f75cb" xmpMM:DocumentID="adobe:docid:photoshop:e72381f3-57f3-d443-a2a9-c45b5b4ac1a8" xmpMM:OriginalDocumentID="xmp.did:aa40acef-ee97-6e42-a032-d944ef89f65e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:aa40acef-ee97-6e42-a032-d944ef89f65e" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:03d57e26-91b7-5440-a88f-df46974f75cb" stEvt:when="2022-09-01T11:02:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>?��  �IDATxڭ��OA ���(�]H$M[z!�48HD��41!R�ME�/0Q�Hś��'�
��@�LC4(>������D�v��Ό��>�-���N�;����o���tclo>�����c�"�eY��t:� GK;�N���x!s���6#��HHmA�P��nǛ=��@�
���D�Sп#	*�u��5�'pr*8����~�� ��lT��qC>��ڰ�+�|^E��6��򅳳�SI?���0�����mn<{}Wp"0}bܞ\����p|�^���G�GI-Ο���z��HR�Uw���\}���BTO^��z��hGpqq�8&���P�^0f1[��J�@�G�I����f��ht�*;>���:&I�\AA>0���f�I�^H���0��!�PRQQ�A��,+�����D�lW���(� ��l�2���Pf8� �fӎ�VBX6O�W۴��t%2��l6Ӆd����`��2���V�
�	��y�5v{��&&h���.\__�[����km�dyy�D"4e��{��Rf�d����߽�����R�8Ք9�jk�Z����=L��-�ب��̀�;=��8�5e�cWm�����3&˱���B!PYY�$)��єy6_p�r��!��2�L�H]����1T#L�jʬ��vi��'C����{X�TOw\�)�����Ӏ���qIt����UD�跑�b0��:�>��a��F�o�?�vtt(����\��A��I    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
�	  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:15+01:00" xmp:MetadataDate="2022-09-01T11:02:15+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:65df7fcf-e4f0-1745-8335-69754b25f309" xmpMM:DocumentID="adobe:docid:photoshop:9b2145bd-a830-e045-a254-fb6668040981" xmpMM:OriginalDocumentID="xmp.did:d3c68f92-932e-984d-8610-1d73a309a547"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d3c68f92-932e-984d-8610-1d73a309a547" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:65df7fcf-e4f0-1745-8335-69754b25f309" stEvt:when="2022-09-01T11:02:15+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�]�B  �IDATxڍ�}lSUƟ�n��v˜u�#1�D`@�Ȃ�1Gɢ�:d�C����2!�(�e����?41�DM�B�`٘ݺ�R��͆h"A�3t#���:�x��j�&o������yn�K8��!�kpp�is�W]shZ����E�� ��n��v�X�h�lE���޼�����E(p�1ʪ�@��L�:my��e䁀��ȏ���s�	�уL�I�mb��e�y<�Ԗ��o�-��� �g�`�O���uuu�����'�>e����-�-	��S��7Nຼ�����|[G����8j���W_z���C#�����ҭ��<t��;�?N)kke[�}��htqJ��R��Q��J�}�Q�{b��m��\�*J����կ��x��ɔ,+β�Rx<���G���Y�1==m^uW����~�/w#c癦���r�������O!<{��g���p��x������o�ָ�˻��Ș j��tA�*-����81�ĩ�Q3oFŞl�&s�r��w}<`��#LU5S�$I&L���߅��J$[gY�F��՟�����Ҫ��� ��P��
�^�	L$�
m�#��Za�J��ޕC�39����L��,�S����<��W��ë�6s0�����9T�,Egt�����Y�0`fh �;��P�!�+߈Y�/\I\�s��A�c�����ŷM��-���SB�J\n�
�/�g3�A�S�b�5�I���X�9�G�_��r�Rm�B_ֲ۰\�U(��n\&!�I��9,����W�v <��Ӹ��� ��²�̰*���&_�
V=�,v�8����h4�u�� �H�r�d���i9�"Vn3Jg��e�6p�h��W�7KPHmRi5������Jh�0��cj���-���2P\{a��ko+D�#��}t�Y�b���vn�3    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:18+01:00" xmp:MetadataDate="2022-09-01T11:02:18+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e9a2bbc4-6b9d-b748-b290-80e6801150a2" xmpMM:DocumentID="adobe:docid:photoshop:e5247389-e03e-804b-b937-37242c86c462" xmpMM:OriginalDocumentID="xmp.did:ac4254a6-7ecf-ef42-b9b8-b23c6b238ffc"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ac4254a6-7ecf-ef42-b9b8-b23c6b238ffc" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e9a2bbc4-6b9d-b748-b290-80e6801150a2" stEvt:when="2022-09-01T11:02:18+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>R�E   �IDATx�c���?��Y��3������G �Y�0Sc�*�31˗��x2�h}�=���C�P�D�ғY)2�p������k�o2;q��i��x J��0f�5Vfpp�9I�59��MRYiIG(6	��LKb%*a@��ˤ�Ȉ3%0L�9��$E����r�"�@\I
FSd ��0y�D���E
AӠ d  ֈF��(�    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:47+01:00" xmp:MetadataDate="2022-09-01T11:02:47+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:da7f1397-745c-9044-8c90-4aebc31c26a4" xmpMM:DocumentID="adobe:docid:photoshop:89924eba-5952-834e-b596-7b986bbf4e12" xmpMM:OriginalDocumentID="xmp.did:0aa08317-5594-cd42-b057-235e4e9adf08"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:0aa08317-5594-cd42-b057-235e4e9adf08" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:da7f1397-745c-9044-8c90-4aebc31c26a4" stEvt:when="2022-09-01T11:02:47+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�r1;   �IDATx�c���?��Y��3������G �Y�0Sc�*�31+�ן�{2�h}�=v��K�P�D��ғ�)2�p���g��7��8���0c��T��@��Kal�0D(I�h�MRT19Ie�%!��D�2Ӓ��J�Ħ ����D�e�ddę�͜Kt�"�@lFu��*U\�l(�aH���M��� ��O���8    IEND�B`� 
BackgroundclWindowNamePaste rightsPngImage.Data

  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:49+01:00" xmp:MetadataDate="2022-09-01T11:02:49+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ec98d2b6-2dae-0347-9ace-568e57646bef" xmpMM:DocumentID="adobe:docid:photoshop:889d205b-3f01-d042-9a6a-6ab3f85584a2" xmpMM:OriginalDocumentID="xmp.did:4415febf-f6c4-d946-b4c9-8186f176322b"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:4415febf-f6c4-d946-b4c9-8186f176322b" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ec98d2b6-2dae-0347-9ace-568e57646bef" stEvt:when="2022-09-01T11:02:49+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�$��  �IDATxڝ��+Q��mV~>(e���D"��XQZ�(ŃMd�$�H��I)���Qh5���$B�Z�Y�3Ύ�1�;�fN��s�����{�D�$ �@��ka$Ɖ���l��"�̢?�R1q��{LWGYn��8�fk0s�����O�_U�����#�$)��b3��U>� ��a�u		�"�1��{�-��`Q�
,f�ń)p��B\l �D�����E~y�z��JL���] �|�t��W�~E�B�{}�����(?JuPO��V{[�rpo�xP�.�8�-�M����0�L�����6N�+Զ{��7���V]�ۧ ��[m�2p{ RZ>����/�;ϫ�Ɔ:�Ř���V#7��{x�MW����F�/0�t/r�jMQ����k��/s(\롷|�g@���~m��(\�
W�쥻��N���-4�p��lᐫA`�9��^l�&&RDZ���o�t��Ku�    IEND�B`�  Leftp  TPngImageListRightsImages144HeightWidth	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:10+01:00" xmp:MetadataDate="2022-09-01T11:02:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:05a047f4-d490-6443-9696-eea015bbb1d5" xmpMM:DocumentID="adobe:docid:photoshop:0d505572-294c-8d4b-b12d-7809f3a4d7c4" xmpMM:OriginalDocumentID="xmp.did:d9ff81b1-dd65-9c47-9f29-780a3c85ff84"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d9ff81b1-dd65-9c47-9f29-780a3c85ff84" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:05a047f4-d490-6443-9696-eea015bbb1d5" stEvt:when="2022-09-01T11:02:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  �IDATxڕ�}leǿ׻��̮�ZVQ@/4FĠ���,�X��2A����h4���A� !��4��m����b� �bT&��]ױ���z�<>w}نe��<��������^�k9J)��8�;<O�AHy��J�B��п�FQ�XSPЍI7���c5(9�j�����I��v�PB>\]�_��gϵ��;ǘ�a� ��*!��+^���gZ[����I����>��J#s�v�
��mv�iuE��⦇�mi?DT�Yg��Hdy~������uOR�t���:���Ғ�_| ���Uxi)��j��
Uݕ����d���c�7ģ��8����gR@}s�L��e3B���#���B�=oA�i�F�ռMe�������(=�+E
e�\.�����q�o�w��� �ظ��}����ʼ�JQw� ^��ȴ�5�w�!�/ͺ��yW�D��a)f�qkj�;�/$t]�v-4zV۽���2��[׭��+j�r}}�)~dY�RkR@��.Q�%�昙���4kBH/�6c��k}�$a�?�x�V���%tt�$J�l��3
H� ���;�mEJ��rc @�5�?���s�7l�=*L �v\`ȱ�H�Eq���-H������B��&I2�1���H?�?��f��C ��΋�9
�g¦E�g����'���u\�?eE���P���=E~�_�5�,� ��`@#� gϵ�5PU�ÞH�6���Ʊ�G�Pak�]̞aA� W�ʂ%��^�� ff��v"R�<��|r��ܒ��nK�6����m�>�흅9���3(���+��܈v^U��.M�?E>�����f��ōC*v�^�_��J{W���4�a�R����݌U;�%�M:@�8`\�~�g��8��~M�����vPA��e.+E������X4A�m�M�G}�)bC�F�_����Ω2�! ��ɾ�9��zwUr@Mm�X�Z��b�L\p��4s>q
��/���N��ۣ&СaW��$5pלJ���p$R��Bp���Wa�)�<r��������r�)"K�P$R�A& NT�����A�v�Y!�s6���R�9�]��T��ރ�ZT;�?,�_�cmG��"�ߡU&����S��PTbb��(#d�-�Y���eu[�0+�K��~��Am]0�&��8�YSl��\tt~�m0%$��{�ߖ�ý �G���P��'�3Q[�%��_Zۄ�>���    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
�	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:13+01:00" xmp:MetadataDate="2022-09-01T11:02:13+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:35ee0ffa-abe8-8445-9ef1-8a089045f471" xmpMM:DocumentID="adobe:docid:photoshop:6132b8cf-07ab-da43-91c0-d89c1c7f8dad" xmpMM:OriginalDocumentID="xmp.did:f75ccada-b4b2-7040-acc4-2f3452e4448c"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:f75ccada-b4b2-7040-acc4-2f3452e4448c" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:35ee0ffa-abe8-8445-9ef1-8a089045f471" stEvt:when="2022-09-01T11:02:13+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  �IDATxڵ�_lE�w��kۣwcP���%�D��\K�-���
�`�bD�
�L�>4��`�PS�R�-m���C�>�))w�&`�ݽ�fv�_/ӊN2w�����3�?3BX���@�H��e^���W�	ވ1�L����=nom��o�i��l ��&B0Pq:	p���N0>�P��?FƮ��'=T����0���qϱ'\��x^�ޟ�H�)�Q�+��!��v�q�K�8�APU���'��������i����F���iH��_ ���1 O��4��drB���>!��HB'�5;ς`|�ꭡ�ZQ]y.�H̬
� �./(�y�����W �L�/����Tc-�G5�C���7{����+]]X�Ų��辘���nb�?�v�gE@gg�\]Sש��qI�A�%Cg}>�?�$���u73�ϯ_ZR���X���pee�!`��۷*�����a͚�Xɜ���ۚ��{��2R*�ң�m%B���ӊ��~�����2�Ȧ����PU�rs`խj�k!`r�E�4?kO(]&T(��j���v�.LLޢhf!(p �D��PUr.@t�b����
u�P,��������aqq�;>���f�x�rY�'Z-���0j��P8d����z/AOw�aoٺ�|t�ׇE�1@���v���q;�P�I�w~�::����?�H$b��H������Q�j��-�f��)�3��/�.���e�Eξmn��� ��,��M?9s2�8w����FYW��5�}Cf�G�.�Lh��2���C<Ѷ�MU��@|�^1��o�IQ�E��u���¶U+E� �oR�����a;EV��~���]�sEp��U��R�CEQ�fNe�$�.�D�ݻ!f��<��Ef��>_�閥���u��($�t�vn9�j���}��^���H~�>ӽ������v!����A���8�    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
�
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:16+01:00" xmp:MetadataDate="2022-09-01T11:02:16+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ce319029-3148-064c-9d86-eaa255a903f4" xmpMM:DocumentID="adobe:docid:photoshop:5efb82e8-7831-ff4b-90f6-b9a0ae42d8f5" xmpMM:OriginalDocumentID="xmp.did:da590269-5f86-da48-b8e8-dca24e9a756f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:da590269-5f86-da48-b8e8-dca24e9a756f" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ce319029-3148-064c-9d86-eaa255a903f4" stEvt:when="2022-09-01T11:02:16+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��,  �IDATxڕ�{lEǿ{�׻����]C���$&`MP��`�(�b���h4���`�5$�@����R�Aci�^[ii��Z5RPQC-Jy��������8�����Q�$s3���g~�ٕcH4I�0��B!�Cq?���PF�SJ���?)H�j��`�&Mh��.��e�(�8��9�F���5�]��v��F�� q� �TsB���V�6m�睝se�����-���'�h����p?���=q�����ֵN��ѵ�����V��?��qc0�4�ɴ���2!��Un\��?55���ˤˌ�
B�ŏ�H�����b��h�f�s����O	hno/P�<O(�:�_Z��T������#\cFܞo��l�p��u����ĩ-2s�ڵWnU%���rۻ�-l~��Mn	���UV�֪��M�Ȋ�<����Ol�� f���j���hT���Ϟ�~����zJ@��NE�#�����󑑑ɟN��3�>>�籘���fHE{��e�)=_������>�99ٶ��D���qc=#�?Bظf>K�w8���X�b������b.Q�q@�%l"�c�	��+Ր�$�ɴ�_��Й���c��7:����,����� �#m8r�(�$Y2�`-��b"/��8��[���$��'UM� ~<�3����M�ȧ֩-Qk����!f�����,�kln��x��B(�y~;D����s)�+�fqq��goEy����/���_/�&B��~�D�D�� �ܫ��$ĭy�fa׽�#͑���%8=�F �@�X��l���1�+lꆖ��#��,.`�/�K}��v{�T� QK4k5f% V���0�^ô�����D��e(�X�W��^�]�au�> �&�[,X܃\�]�o@4�"<�o-�Ɯ�Ÿ�������qp�M�{lq*<�'�����D����%;y��R��,ŋm[0;�ns�e�^��������@�I��!����!6��* e�;� �d�/n�����S)N_����@0���mI���GUU�x�M�U �9҃�X��D�]�L^A�q!�[�83X��n�&� �1��6M�+�0���[���_y�f�1�J�B��[P�\"2�O*�+�x���tZ�9˟���L�������K\��E���c8a�/<�j�>�    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
7  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:19+01:00" xmp:MetadataDate="2022-09-01T11:02:19+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f0f547b5-21de-b240-8075-d653261399a4" xmpMM:DocumentID="adobe:docid:photoshop:8caa230a-947e-f144-9663-a8ea5172874b" xmpMM:OriginalDocumentID="xmp.did:4dfea257-8368-1d45-89b3-ca52ddae4d2c"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:4dfea257-8368-1d45-89b3-ca52ddae4d2c" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f0f547b5-21de-b240-8075-d653261399a4" stEvt:when="2022-09-01T11:02:19+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  IDATx�c���?��Y��3��
�ӓ�0� @f3�,HI�ũp���,,,_~���I�%$Y�����}��,!����W�I��$�����dV�Y��B���`J `�@�XY�1;q
N��A�Լ���$	3��فa��DY��W�Z �N�c���3���	Z��W�Ғ�� Ƈ��Լ����J�� #5�-`$)Qd1�ȶ���`�a�6s.ə�,��t�l��+ȩ�*� r^���/����,����
�-@�+�3m:�,  �!��(ό\    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:47+01:00" xmp:MetadataDate="2022-09-01T11:02:47+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:028ed0ca-db2d-b446-b46b-d7506905e41a" xmpMM:DocumentID="adobe:docid:photoshop:b414145a-2a3e-414f-86d6-295fc78c6358" xmpMM:OriginalDocumentID="xmp.did:9dadd350-edd7-3d43-b2c4-6ded0d027b9e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:9dadd350-edd7-3d43-b2c4-6ded0d027b9e" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:028ed0ca-db2d-b446-b46b-d7506905e41a" stEvt:when="2022-09-01T11:02:47+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�K��   �IDATx�c���?��Y��3��
�ӓ�0� @f3�,HI�ũp���l��_���A�%$Y�����s�^�,!����W�I��$�����df�Y��B���`J `��]��p��)�������:����A7���
Q���,@�+YiIG��,�I�+�iI��X`�h#I��"��D����ô�sIΌdY�/�P�|y�f`KiT���O�8���dY@��P �  �������M    IEND�B`� 
BackgroundclWindowNamePaste rightsPngImage.Data
}  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:50+01:00" xmp:MetadataDate="2022-09-01T11:02:50+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:5e812b52-cf2a-6148-935f-ff86be43b13c" xmpMM:DocumentID="adobe:docid:photoshop:9a416c63-fa66-164d-8373-443e53795f0b" xmpMM:OriginalDocumentID="xmp.did:2235ab72-75fb-4846-91e7-912edaab2d19"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:2235ab72-75fb-4846-91e7-912edaab2d19" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:5e812b52-cf2a-6148-935f-ff86be43b13c" stEvt:when="2022-09-01T11:02:50+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?><���  ZIDATx�c���?0222`����r-b�����̯�b���<c ��f$d��=��3�U�`d`қ�\��Sł_�$M���R<��3��p0�c��?��������D� %��@�H��������`����d��������c����#�(�����@� U���?/�1��򈁛h#�p���'��{�}\��Cr����X��s�.N� ��7�8ЂWx-�r~�b`x��x�X@ �0�C� K�	���� �˂� �c� ����ś$Aq���itzn�2�mF� ��7d�2�$��`���,��?�������Â#M�} 7�[�����m��~�v��H9�b���q ·[ ���5���{�����=+-�܂C��/��	�;��._�����c"C� ����̴$f��P-@����� ���0�-�W�x��
n���P,�[����@�B��ɏ�)���
H2E�\~�A�v�c�d˞hR�e���g��`{	$��
��:�`[1�| ���.�>�R�x	���D��)�`u#�~A\>��}A��P �  �d�)vH    IEND�B`�  Leftx  TPngImageListRightsImages192Height Width 	PngImages
BackgroundclWindowName'No rights-preset on permissions controlPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:11+01:00" xmp:MetadataDate="2022-09-01T11:02:11+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b1cae5af-18fa-6c42-aae1-7c7f937c2bee" xmpMM:DocumentID="adobe:docid:photoshop:cc4155c3-b9cb-fb4b-86f8-a28545dc7f23" xmpMM:OriginalDocumentID="xmp.did:a9d6e70b-6ba5-3241-812a-1d9ace758465"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:a9d6e70b-6ba5-3241-812a-1d9ace758465" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b1cae5af-18fa-6c42-aae1-7c7f937c2bee" stEvt:when="2022-09-01T11:02:11+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>K�QB  �IDATx�͗}Lg�WJ��D@���n&&.�I�f����!/
3��6gܖmYb�ɲ?�����6�w���D�������"P{�]�=�W���:4۞�����<���{{R
!���� E�����(}�����ݻw�$/I@���DEJ���!�*�X�C뵓�N|� ����(QwLDh,���[�+槥��|f ��/�R�+��o���.A�2׭=�� uuMs��`;S�8�p�@4jx�ɋ������� ���EK�!�S�c�"�
׬I�%�UUW�1d'΁� ��2�����i5�V�Hܺ:e���*���a�C~��,'+�v\ �����}�*Υ�R�n�D啧*��� ���fg������,%�pv�OM]~},����d��5�J���y�YI��P[�bq��Gm��5���4)�"���8�6�@�E+Rg��U˃j�ߝ(GJ����٣��܅:�N���)A|[\���͜p�Ƕo\.gn&d����`t�2:::�<�4MK^��[A\i��/
�'(vri���3�; ��F .{m1@��n�2 �9 @~�nmwC%���H��uۆ� C�X�*U1�]�]|�sV��r3R����8�S�O˵6���!v��3_�.���6�?�k��t,c�1NMv?�q��zM����1 ��\�?���ﷂ�9tw���1&�<H<!y@����0��+3Ѱ�<+����v��:M �	��8>>���Қ���p��~��~�QO�`�t�l,��������a�90�(��;����L׃?X�ŵ�Y�JM���U�'$�N� ��n���Ab?u�؛d Cw̈����M<џ���T\ a}w��@��,��D<�8M u�K^HHP d�Kk�m�G/���������)|]m;� �^�Ƒ5a����hl]�������Zgj."��	�	�mu���>��b_��l�۽���="
�@/р�H�{�.�Z|T��gϫr i �嗕�N�K��G�������=yo��ǿ��j�QN�>�|�� �2�}qI�pS�D�N���'�d�~���q��� *O�QH!HT5"����m+���rX~�C Zva��0-�ြw�$��9��j����H9���#���8��m&�cHG�.�p�o��ϱjQCh�V�B��\HL
��R*�����m�2	�p���<:Wn'룿�J�C�x�e9nB�DY�_'LLJSHX��ı�#/������"��M�.{��Al�>�b��FN
a���@h�V"A|I8��|# !G>��i��c �YG������!�G�-V:T�0�L��=^�݊O��9������.�᡾������G!�B00-��N�%+��& *�L(6�I�C�ք�dW�����q�����j�B�{<\Z`�rӆ*����0�h֪    IEND�B`� 
BackgroundclWindowNameDefault rights-presetPngImage.Data
'
  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:14+01:00" xmp:MetadataDate="2022-09-01T11:02:14+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:bf3f4354-ed1c-fd4e-8bcd-90c671ae8e4c" xmpMM:DocumentID="adobe:docid:photoshop:2e158c41-5867-644b-ba03-36fd0913e7cd" xmpMM:OriginalDocumentID="xmp.did:1e743dfa-4102-434d-9cda-6886d1496e52"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:1e743dfa-4102-434d-9cda-6886d1496e52" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:bf3f4354-ed1c-fd4e-8bcd-90c671ae8e4c" stEvt:when="2022-09-01T11:02:14+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��R  IDATx�͖�OA�gkb�h�z�,}�LLHP4�T��J�Riim$Q�z�1!���S
EBQT��P=@|�DL��4��83��ζ�2T�nӝ��o����=�B��K�/A�����H������kj-���Y�u{Y-��!X
!�@���QD���o^���v��	Pw"�	,����h���m��@��3� tA,�*]���oU��(Bg]�����lF:0��V����wH`�Ǝ���?�������KJ��DE�8�ß���:A���M �8�c��2^_W]�3���H%��"�G*���ZA��n�VWU;���v '�����������j�Y��PwH��F�2N��q9=�D�>bo��Gw��V>����s;��IW���u9�9<����d�~���_�贴t�^�^���dn�ކkr�{���m�(�*�w�u �d���rx�8�؀�o�r�U�������[�^\L�$���<���ԔXB���ܶ���`�N}(*� �vRj��>� �>%(����];.����-� �9@�w5 n�D��ղ�`�Y���`(T�Zk���Jяj�}�� "C#Y R�!=���)��N��b@�Ƕ���+ �ժɘ��(�|�"͘c�O��%%��&�q��c���<�dҏ U+#c��07;K�׭[n��.	PU����2�h4f����a03�����[� ���8`穩����=A���&�jb�<99	Μ>E�Ϟ;�m̩��sf8��| =11�4 ��s:j�}[�C���N�8k�� ��<D�i���YG�mAe�,H<K��4�s���e �Lꢓ;�t��_i�� ���������Z JĘ��Gr� �1�h��Fl1�MY�2+��.�V�O�>O=��`HU	Mf�bZ;��V2�|�cyI�@{���O
 ML��# )W"��k�̂޾��s�����ᓼ��(k���S �+?U��i����/x� tŘu    IEND�B`� 
BackgroundclWindowNameAll rights-presetPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:17+01:00" xmp:MetadataDate="2022-09-01T11:02:17+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:98c9ccf1-a9d9-4049-bdae-58b68d7ee6e9" xmpMM:DocumentID="adobe:docid:photoshop:f53c22ba-071f-1541-b51f-45fded1f96f8" xmpMM:OriginalDocumentID="xmp.did:6658f49f-d6e3-0046-a110-e8dc60d61ffc"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:6658f49f-d6e3-0046-a110-e8dc60d61ffc" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:98c9ccf1-a9d9-4049-bdae-58b68d7ee6e9" stEvt:when="2022-09-01T11:02:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  �IDATx�͗{LGǿ�wp �@�Fl�E�&hC�1%�(�'&�� ���Q������-M�&ڤ�6�i��7o*�C@��Z����r���y�;���{�Rj�.agٝ������QJ�_^����!-����ƌ�ۿ����ύ�Mh�d>!t���=D��$��҅B6��p�������Jg2A0q��>7Q�d,[�����W��s�s�����Ҩ����*�$9i�ғ����6��8��(�n6"?�X�I_t�ׇ �|��������L0��⛤y��3A4�X� iX��,z� յK�x���HɆ%�q?�m�WP������S�S�+�P~���������q��(7�x�H�r��:�pZJr�� *�[Y�_s$��h�~Q�` ǎ��P����J������a����a�~��v����yMg�޼�c�8�,.�͒1}��Q�();C�3;a�!��CGs�#�ڌ���8u���'�R}�� �� _�n���|����jIg�D�$44t(��\���J0	�N�?fC8w��>�Np�SJK~P��tv>�\��mnH 5��S�� �; p����NK+���o��f���3S��ĕ�3*��=��lu��Ӧ�zX�f�@�Qp�+\�n��������M�Qk'�K9���e\ۜ�>� �յ� ���|�p{/��Qӊa6H9,oK]��ˢ
s��&��|��h��
�:��$a �<�����������3oS0�c�! ��C�]\� �:n�.�Ԫ����gLU(-�r+?	 �i� =m5�&s�����1>�_�ϊK�ۧ�㍱��˫p��E����/J���%/��9 �Kk6�_��/-0aR�!ԫ���l�8����/E��g���#=]�>U�%e���EXx���� ZZZ���O��!ƿ��?�%�)���㛨�����o����oKLK���*@��R��* ���+��� p���Ҙ8��C>D���7Ƃ{YB>��UO�¢S�y��*9I�#  4`6f�Q|ol�SL�{;��sZY�����T�^ �p�B��t��mڸ��4�Z�u�?"&x%n���y)��~�ccQ��a�k��������Q��j ΎȞK;��M�R�M$�;�E��cw�]�^�o[��x�<�o�n���$��;N�K���vOt�:p�eFEZ�2������,���+�U"��+C����{t�����= �㩻��&���҈��>�Qco'���DI<Gr��z�ވ6{iDG��(��$t8N>O ��#��#<�ށ�e��uD�s���{+�c�V\x���dN�u� n ��w��O���N���>���k�i�;�f��46掂�q͠��P�9U���Fj��l�x�`y?L�L����_|��̟&    IEND�B`� 
BackgroundclWindowNameCopy rights-permissions as textPngImage.Data
[  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:17+01:00" xmp:ModifyDate="2022-09-01T11:02:20+01:00" xmp:MetadataDate="2022-09-01T11:02:20+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f1541377-eda2-9047-94b4-013022ed231f" xmpMM:DocumentID="adobe:docid:photoshop:ae4447a8-a9c1-9546-b293-71aa366f0e75" xmpMM:OriginalDocumentID="xmp.did:c0ca06a3-2ffa-4b44-ba5a-6c25b74d12da"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c0ca06a3-2ffa-4b44-ba5a-6c25b74d12da" stEvt:when="2022-06-27T15:59:17+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f1541377-eda2-9047-94b4-013022ed231f" stEvt:when="2022-09-01T11:02:20+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>+YŖ  8IDATx����KSa�����ηj�(1Tz�1�2���Pj(��c���A *˵2�%VVC��m�����΋��6�ǝs|�n��=p���<��+$�I�3Bp�����=624���C��9pC׀{�S�X,�U�0���v^�?�h
��]��f
�����utd��H ,�90�?+��:4అ�03�CMU%B�먫ub{{�<�Y�����
�n,-9�Ɔz�lV�Bkp8�q���0�VX� �<dӲ�zc3B����:�SӆZ�#F��Y��^�u<G`�Z�\Xx������`�����/D�=sד�9TWV�ShU7��"����:���dY�`3���e$R��	Bꀜ��@�=����GȒ��g�!I��_��{��=nZ����UX��O��{��ۅ����Q�[���
˷��(�BN���%�nR� Vai���p:Obi�=:��P\\��*,Q�+P���O|ݍ��@�y҅���	�����Q�<��f�� ҅u��Zj���cx���(/�8��X�
0. ӻ����z&r�&�)    IEND�B`� 
BackgroundclWindowName Copy rights-permissions as octalPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:48+01:00" xmp:MetadataDate="2022-09-01T11:02:48+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:97e1dd6f-4b03-0143-846d-1ea8a9d02ebf" xmpMM:DocumentID="adobe:docid:photoshop:454835e8-b3b8-9e4e-b1d6-3ecbb4d9c273" xmpMM:OriginalDocumentID="xmp.did:72e32afa-ca30-3f4a-a59d-0617ca72282c"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:72e32afa-ca30-3f4a-a59d-0617ca72282c" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:97e1dd6f-4b03-0143-846d-1ea8a9d02ebf" stEvt:when="2022-09-01T11:02:48+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>: ��  �IDATx����Oq��������~Y��責f�i��_K�.�j���zVR�[ITk�@:5�?X�Px4:ny�u'�;��Z�'w�}w��}��yS�|[Y�:����b$?��mW�{R6���� �/�'z��;��T*S�\�,!�j1��&	!����RLB6@�� d�Tn���� �P���4 �N��h�x4M��^�V]�����C�\�hԨ��Cly^�SX�'P]]�6X�����F|�p�4
����������c7R��( _`	�i�x(���-�LL"����v,Ŗ��xE�K�bl���Yt�,܂��)�~�Cg�Y�/����� /��@8G���R <�����V��|���ϝEQ�P�h��{� �b ܸ�1�.��4��C<��g��M�����?��=��h�{U�*@�فյ5<�
+�xy$/ 	��J�$ iI�V�e�3�,��n�ٵu{w�O}��vc�(�<�4�d<A&������ 	��!LMπb:�[�M� 	�dr����q���� 	,�Ǉ��*��/���Ď�l ��Z\������(��8�m���J� ���fn$_�A�M�榃��ֿ�����lU�4���=    IEND�B`� 
BackgroundclWindowNamePaste rightsPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:50+01:00" xmp:MetadataDate="2022-09-01T11:02:50+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:2f5b12d6-947b-b041-ba3c-933440bb754b" xmpMM:DocumentID="adobe:docid:photoshop:ba0be574-3911-f142-bd60-3dda6723a7a1" xmpMM:OriginalDocumentID="xmp.did:c2e157e7-6f02-6749-8eeb-b77b8fe8423b"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c2e157e7-6f02-6749-8eeb-b77b8fe8423b" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:2f5b12d6-947b-b041-ba3c-933440bb754b" stEvt:when="2022-09-01T11:02:50+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��j  zIDATx�c���?0222�WW1��H5312D�����_x���F�0�_$ ;Iq���R�@%(�1��`w}^I��#���F	���X��:u<cu}&MS��*��������"�ג����L,G�������{���[9�D�' ŋ���L�(�����M����j��u�l��*6��@&@�p��ӭ��?c�H�03�C3#�����{�Fu ��Q� ���9qQ r�� B�h�v2 џ�)��W���  �� ����؄Թw�㭄pUj.qAL��$�t14�&��Z\\�&=�!%1�(̙������Ͽ,����G:�h3a\�!����w�����O�#p:�H~��M9� R���kG�t��F��%O�@ �YiIG�:�P���� Y���������Ċ��	;��"�!�+T���
��p�E�]%�B [�t��Z���L��WC��Uh{�	;��*C`Oa<T�a�$�G�4�]����A��YN�O4i;��O�h�K	;��6C`k1j���C`Ka�Хal.`<l�Y�K�/�h� B}C�6s��� �  ��߃��:    IEND�B`�  Left�       TPF0�TScpCommanderFormScpCommanderFormLeft� Top HelpType	htKeywordHelpKeywordui_commanderCaptionScpCommanderFormClientHeight�ClientWidth�
TextHeight � 	TSplitterSplitterLeft�Top� WidthHeight!CursorcrSizeWEHintj   |Dra för att ändra proportioner på filpaneler. Dubbelklicka för att bredden på filpanelerna ska lika.ResizeStylersUpdateOnCanResizeSplitterCanResizeOnMovedSplitterMoved  �	TSplitterQueueSplitterTopWidth�  �TTBXDockTopDockWidth�Height� OnContextPopupDockContextPopup TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	OptionstboNoAutoHinttboShowHint 
ShrinkModetbsmWrapStretch	TabOrder TTBXSubmenuItemLocalMenuButtonCaption&LocalXHelpKeywordui_commander_menu#local TTBXItemTBXItem1Action*NonVisualDataModule.LocalChangePathAction2  TTBXSeparatorItemTBXSeparatorItem1  TTBXSubmenuItemTBXSubmenuItem2Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItemTBXItem2Action&NonVisualDataModule.LocalOpenDirAction  TTBXItemTBXItem3Action/NonVisualDataModule.LocalExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem2  TTBXItemTBXItem4Action(NonVisualDataModule.LocalParentDirAction  TTBXItemTBXItem5Action&NonVisualDataModule.LocalRootDirAction  TTBXItemTBXItem6Action&NonVisualDataModule.LocalHomeDirAction  TTBXItem
TBXItem262Action'NonVisualDataModule.LocalOtherDirAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXItemTBXItem7Action#NonVisualDataModule.LocalBackAction  TTBXItemTBXItem8Action&NonVisualDataModule.LocalForwardAction   TTBXItemTBXItem9Action&NonVisualDataModule.LocalRefreshAction  TTBXItem	TBXItem10Action+NonVisualDataModule.LocalAddBookmarkAction2  TTBXItem	TBXItem11Action/NonVisualDataModule.LocalPathToClipboardAction2  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemTBXSubmenuItem17Caption&VyHelpKeywordui_file_panel#view_styleHint   Ändra stil för katalogvy TTBXItem
TBXItem270Action%NonVisualDataModule.LocalReportAction  TTBXSeparatorItemTBXSeparatorItem76  TTBXItem
TBXItem271Action(NonVisualDataModule.LocalThumbnailAction   TTBXSubmenuItemTBXSubmenuItem3Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i lokal panel TTBXItem	TBXItem12Action-NonVisualDataModule.LocalSortAscendingAction2  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem13Action*NonVisualDataModule.LocalSortByNameAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem14Action)NonVisualDataModule.LocalSortByExtAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem17Action*NonVisualDataModule.LocalSortBySizeAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem15Action*NonVisualDataModule.LocalSortByTypeAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem16Action-NonVisualDataModule.LocalSortByChangedAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem18Action*NonVisualDataModule.LocalSortByAttrAction2
GroupIndex	RadioItem	   TTBXSubmenuItemLocalColumnsSubmenuItemCaption	&KolumnerHelpKeywordui_file_panel#selecting_columns TTBXItem	TBXItem19Action2NonVisualDataModule.ShowHideLocalNameColumnAction2  TTBXItem	TBXItem20Action2NonVisualDataModule.ShowHideLocalSizeColumnAction2  TTBXItem	TBXItem21Action2NonVisualDataModule.ShowHideLocalTypeColumnAction2  TTBXItem	TBXItem22Action5NonVisualDataModule.ShowHideLocalChangedColumnAction2  TTBXItem	TBXItem23Action2NonVisualDataModule.ShowHideLocalAttrColumnAction2  TTBXSeparatorItemTBXSeparatorItem72  TTBXItem
TBXItem263Action.NonVisualDataModule.AutoSizeLocalColumnsAction  TTBXItem
TBXItem265Action1NonVisualDataModule.ResetLayoutLocalColumnsAction   TTBXItem
TBXItem221Action%NonVisualDataModule.LocalFilterAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_commander_menu#markHint   Kommandon för markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXSeparatorItemTBXSeparatorItem60  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction  TTBXSeparatorItemTBXSeparatorItem61  TTBXItem
TBXItem212Action'NonVisualDataModule.SelectSameExtAction  TTBXItem
TBXItem213Action)NonVisualDataModule.UnselectSameExtAction   TTBXSubmenuItemTBXSubmenuItem5Caption&FilerHelpKeywordui_commander_menu#filesHint   Kommandon för filoperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem	TBXItem28Action!NonVisualDataModule.NewFileAction  TTBXItem	TBXItem24Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXSubmenuItem	TBXItem26Action%NonVisualDataModule.CurrentEditActionDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem	TBXItem29Action,NonVisualDataModule.CurrentAddEditLinkAction  TTBXSeparatorItemTBXSeparatorItem7  TTBXSubmenuItemCurrentCopyItemAction$NonVisualDataModule.RemoteCopyActionDropdownCombo	 TTBXItemCurrentCopyNonQueueItemAction,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItemCurrentCopyQueueItemAction)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem51  TTBXItemCurrentMoveItemAction$NonVisualDataModule.RemoteMoveAction   TTBXItemCurrentCopyToItemAction&NonVisualDataModule.RemoteCopyToAction  TTBXItemCurrentMoveToItemAction&NonVisualDataModule.RemoteMoveToAction  TTBXItem	TBXItem34Action'NonVisualDataModule.CurrentDeleteAction  TTBXItem	TBXItem35Action'NonVisualDataModule.CurrentRenameAction  TTBXSeparatorItemTBXSeparatorItem62  TTBXItem
TBXItem163Action1NonVisualDataModule.CurrentCopyToClipboardAction2  TTBXItem	TBXItem36Action NonVisualDataModule.PasteAction3  TTBXSeparatorItemTBXSeparatorItem8  TTBXSubmenuItemCustomCommandsMenuAction,NonVisualDataModule.CustomCommandsFileAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem37Action/NonVisualDataModule.FileListToCommandLineAction  TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action*NonVisualDataModule.FileGenerateUrlAction2   TTBXSubmenuItemTBXSubmenuItem25Caption	   &LåsningHint   Hantera fillås TTBXItem
TBXItem214ActionNonVisualDataModule.LockAction  TTBXItem
TBXItem216Action NonVisualDataModule.UnlockAction   TTBXSeparatorItemTBXSeparatorItem9  TTBXItem	TBXItem41Action+NonVisualDataModule.CurrentPropertiesAction  TTBXItem
TBXItem239Action1NonVisualDataModule.CalculateDirectorySizesAction   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_commander_menu#commandsHintAndra kommandon TTBXItem	TBXItem42Action-NonVisualDataModule.CompareDirectoriesAction2  TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItem	TBXItem45Action.NonVisualDataModule.SynchronizeBrowsingAction2  TTBXItem
TBXItem210Action*NonVisualDataModule.RemoteFindFilesAction2  TTBXSubmenuItemQueueSubmenuItemCaption   K&öHelpKeywordui_queue#manageHint   Kommandon för kölistaOnPopupQueueSubmenuItemPopup TTBXItemQueueEnableItem2Action%NonVisualDataModule.QueueEnableAction  TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#manageHint&   Administrationskommandon för kömassa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction  TTBXItem
TBXItem142Action(NonVisualDataModule.QueueDeleteAllAction  TTBXSeparatorItemTBXSeparatorItem39  TTBXItem
TBXItem134Action,NonVisualDataModule.QueueDeleteAllDoneAction    TTBXSubmenuItemTBXSubmenuItem28Action/NonVisualDataModule.CustomCommandsNonFileAction  TTBXSeparatorItemTBXSeparatorItem13  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction  TTBXSeparatorItemTBXSeparatorItem15  TTBXItem	TBXItem58Action+NonVisualDataModule.CloseApplicationAction2   TTBXSubmenuItemTBXSubmenuItem29Caption&FlikarHelpKeywordui_commander_menu#tabsHintTabkommandon TTBXSubmenuItemTBXSubmenuItem30Action NonVisualDataModule.NewTabActionDropdownCombo	 TTBXItem	TBXItem33Action&NonVisualDataModule.NewRemoteTabAction  TTBXItem	TBXItem31Action%NonVisualDataModule.NewLocalTabAction  TTBXSeparatorItemTBXSeparatorItem67  TTBXItem
TBXItem232Action/NonVisualDataModule.DefaultToNewRemoteTabAction   TTBXItem
TBXItem115Action"NonVisualDataModule.CloseTabAction  TTBXItem
TBXItem218Action&NonVisualDataModule.DuplicateTabAction  TTBXItem
TBXItem127Action#NonVisualDataModule.RenameTabAction  TTBXSeparatorItemTBXSeparatorItem53  TTBXColorItemColorMenuItemAction$NonVisualDataModule.ColorMenuAction2ColorclNone  TTBXSeparatorItemTBXSeparatorItem69  TTBXItem
TBXItem252Action+NonVisualDataModule.DisconnectSessionAction  TTBXItem
TBXItem253Action*NonVisualDataModule.ReconnectSessionAction  TTBXItem
TBXItem114Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem50  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem
TBXItem135Action-NonVisualDataModule.SessionGenerateUrlAction2  TTBXItem
TBXItem227Action(NonVisualDataModule.ChangePasswordAction  TTBXItem	TBXItem76Action*NonVisualDataModule.PrivateKeyUploadAction  TTBXSeparatorItemTBXSeparatorItem29  TTBXSubmenuItemTBXSubmenuItem21Action$NonVisualDataModule.OpenedTabsAction  TTBXSubmenuItemTBXSubmenuItem231Action$NonVisualDataModule.WorkspacesAction  TTBXItem
TBXItem230Action'NonVisualDataModule.SaveWorkspaceAction  TTBXSeparatorItemTBXSeparatorItem23  TTBXSubmenuItemTBXSubmenuItem20Action(NonVisualDataModule.SavedSessionsAction2   TTBXSubmenuItemTBXSubmenuItem9Caption&AlternativHelpKeywordui_commander_menu#optionsHint)   Ändra layout/inställningar för program TTBXSubmenuItemTBXSubmenuItem10Caption   &VerktygsfältHelpKeywordui_toolbarsHint   Visa/dölj verktygsfält TTBXItem	TBXItem64Action/NonVisualDataModule.CommanderCommandsBandAction  TTBXItem	TBXItem60Action/NonVisualDataModule.CommanderSessionBandAction2  TTBXItem	TBXItem62Action2NonVisualDataModule.CommanderPreferencesBandAction  TTBXItem	TBXItem63Action+NonVisualDataModule.CommanderSortBandAction  TTBXItem
TBXItem186Action.NonVisualDataModule.CommanderUpdatesBandAction  TTBXItem
TBXItem188Action/NonVisualDataModule.CommanderTransferBandAction  TTBXItem
TBXItem215Action5NonVisualDataModule.CommanderCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem38  TTBXItem	TBXItem74Action"NonVisualDataModule.ToolBar2Action  TTBXSeparatorItemTBXSeparatorItem47  TTBXItem
TBXItem191Action&NonVisualDataModule.LockToolbarsAction  TTBXItem
TBXItem133Action.NonVisualDataModule.SelectiveToolbarTextAction  TTBXSubmenuItem
TBXItem272Action)NonVisualDataModule.ToolbarIconSizeAction TTBXItem
TBXItem273Action/NonVisualDataModule.ToolbarIconSizeNormalAction	RadioItem	  TTBXItem
TBXItem274Action.NonVisualDataModule.ToolbarIconSizeLargeAction	RadioItem	  TTBXItem
TBXItem275Action2NonVisualDataModule.ToolbarIconSizeVeryLargeAction	RadioItem	    TTBXSubmenuItemTBXSubmenuItem11Action-NonVisualDataModule.CommanderLocalPanelAction TTBXItem	TBXItem65Action4NonVisualDataModule.CommanderLocalHistoryBandAction2  TTBXItem	TBXItem66Action7NonVisualDataModule.CommanderLocalNavigationBandAction2  TTBXItem	TBXItem59Action1NonVisualDataModule.CommanderLocalFileBandAction2  TTBXItem	TBXItem61Action6NonVisualDataModule.CommanderLocalSelectionBandAction2  TTBXSeparatorItemTBXSeparatorItem16  TTBXItem	TBXItem67Action#NonVisualDataModule.LocalTreeAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXItem	TBXItem68Action)NonVisualDataModule.LocalStatusBarAction2   TTBXSubmenuItemTBXSubmenuItem12Action.NonVisualDataModule.CommanderRemotePanelAction TTBXItem	TBXItem69Action5NonVisualDataModule.CommanderRemoteHistoryBandAction2  TTBXItem	TBXItem70Action8NonVisualDataModule.CommanderRemoteNavigationBandAction2  TTBXItem
TBXItem136Action2NonVisualDataModule.CommanderRemoteFileBandAction2  TTBXItem
TBXItem131Action7NonVisualDataModule.CommanderRemoteSelectionBandAction2  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem19  TTBXItem	TBXItem72Action*NonVisualDataModule.RemoteStatusBarAction2   TTBXSeparatorItemTBXSeparatorItem20  TTBXItemSessionsTabs3Action'NonVisualDataModule.SessionsTabsAction2  TTBXItem	TBXItem73Action*NonVisualDataModule.CommandLinePanelAction  TTBXItem	TBXItem75Action#NonVisualDataModule.StatusBarAction  TTBXSubmenuItemTBXSubmenuItem14Caption   K&öHelpKeywordui_queueHint   Konfigurera kölista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXItem
TBXItem255Action'NonVisualDataModule.QueueFileListAction  TTBXSeparatorItemTBXSeparatorItem74  TTBXItem
TBXItem267Action1NonVisualDataModule.QueueResetLayoutColumnsAction  TTBXSeparatorItemTBXSeparatorItem22  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action3NonVisualDataModule.QueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem141Action0NonVisualDataModule.QueueSuspendOnceEmptyAction2  TTBXItem
TBXItem224Action1NonVisualDataModule.QueueShutDownOnceEmptyAction2	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXSeparatorItemTBXSeparatorItem49  TTBXItem	TBXItem82Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemRemoteMenuButtonCaption&RemoteXHelpKeywordui_commander_menu#remote TTBXItem	TBXItem83Action+NonVisualDataModule.RemoteChangePathAction2  TTBXSeparatorItemTBXSeparatorItem24  TTBXSubmenuItemTBXSubmenuItem15Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXItem
TBXItem257Action0NonVisualDataModule.RemoteExploreDirectoryAction  TTBXSeparatorItemTBXSeparatorItem25  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem
TBXItem261Action(NonVisualDataModule.RemoteOtherDirAction  TTBXSeparatorItemTBXSeparatorItem26  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem90Action'NonVisualDataModule.RemoteRefreshAction  TTBXItem	TBXItem91Action,NonVisualDataModule.RemoteAddBookmarkAction2  TTBXItem	TBXItem92Action0NonVisualDataModule.RemotePathToClipboardAction2  TTBXSeparatorItemTBXSeparatorItem27  TTBXSubmenuItemTBXSubmenuItem19Caption&VyHelpKeywordui_file_panel#view_styleHint   Ändra stil för katalogvy TTBXItem
TBXItem276Action&NonVisualDataModule.RemoteReportAction  TTBXSeparatorItemTBXSeparatorItem77  TTBXItem
TBXItem277Action)NonVisualDataModule.RemoteThumbnailAction   TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i fjärrpanel TTBXItem	TBXItem93Action.NonVisualDataModule.RemoteSortAscendingAction2  TTBXSeparatorItemTBXSeparatorItem28  TTBXItem	TBXItem94Action+NonVisualDataModule.RemoteSortByNameAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem95Action*NonVisualDataModule.RemoteSortByExtAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem97Action+NonVisualDataModule.RemoteSortBySizeAction2
GroupIndex	RadioItem	  TTBXItem
TBXItem193Action+NonVisualDataModule.RemoteSortByTypeAction2	RadioItem	  TTBXItem	TBXItem96Action.NonVisualDataModule.RemoteSortByChangedAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem98Action-NonVisualDataModule.RemoteSortByRightsAction2
GroupIndex	RadioItem	  TTBXItem	TBXItem99Action,NonVisualDataModule.RemoteSortByOwnerAction2
GroupIndex	RadioItem	  TTBXItem
TBXItem100Action,NonVisualDataModule.RemoteSortByGroupAction2
GroupIndex	RadioItem	   TTBXSubmenuItemRemoteColumnsSubmenuItemCaption	&KolumnerHelpKeywordui_file_panel#selecting_columns TTBXItem
TBXItem101Action3NonVisualDataModule.ShowHideRemoteNameColumnAction2  TTBXItem
TBXItem102Action3NonVisualDataModule.ShowHideRemoteSizeColumnAction2  TTBXItem
TBXItem192Action3NonVisualDataModule.ShowHideRemoteTypeColumnAction2  TTBXItem
TBXItem103Action6NonVisualDataModule.ShowHideRemoteChangedColumnAction2  TTBXItem
TBXItem104Action5NonVisualDataModule.ShowHideRemoteRightsColumnAction2  TTBXItem
TBXItem105Action4NonVisualDataModule.ShowHideRemoteOwnerColumnAction2  TTBXItem
TBXItem106Action4NonVisualDataModule.ShowHideRemoteGroupColumnAction2  TTBXItem
TBXItem179Action9NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction2  TTBXSeparatorItemTBXSeparatorItem73  TTBXItem
TBXItem264Action/NonVisualDataModule.AutoSizeRemoteColumnsAction  TTBXItem
TBXItem266Action2NonVisualDataModule.ResetLayoutRemoteColumnsAction   TTBXItem
TBXItem220Action&NonVisualDataModule.RemoteFilterAction   TTBXSubmenuItemTBXSubmenuItem22Caption   &HjälpHelpKeywordui_commander_menu#helpHint   Hjälp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXItem
TBXItem217ActionNonVisualDataModule.TipsAction  TTBXSeparatorItemTBXSeparatorItem30  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarPreferencesToolbarLeft Top3Caption   InställningarDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem65  TTBXItem
TBXItem256Action'NonVisualDataModule.QueueFileListAction    TTBXToolbarSessionToolbar2Left TopCaptionSessioner och flikarDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder  TTBXSubmenuItemTBXSubmenuItem31Action NonVisualDataModule.NewTabActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem231Action&NonVisualDataModule.NewRemoteTabAction  TTBXItem
TBXItem123Action%NonVisualDataModule.NewLocalTabAction  TTBXSeparatorItemTBXSeparatorItem68  TTBXItem
TBXItem238Action/NonVisualDataModule.DefaultToNewRemoteTabAction   TTBXItem
TBXItem125Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem66  TTBXItem
TBXItem219Action&NonVisualDataModule.DuplicateTabAction  TTBXItem
TBXItem124Action"NonVisualDataModule.CloseTabAction  TTBXSeparatorItemTBXSeparatorItem34  TTBXSubmenuItemTBXSubmenuItem23Action(NonVisualDataModule.SavedSessionsAction2DisplayModenbdmImageAndTextOptionstboDropdownArrow    TTBXToolbarSortToolbarLeft TopMCaptionSorteraDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem148Action,NonVisualDataModule.CurrentSortByTypeAction2  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarCommandsToolbarLeft TopgCaption	KommandonDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem154Action-NonVisualDataModule.CompareDirectoriesAction2  TTBXItem
TBXItem155Action%NonVisualDataModule.SynchronizeAction  TTBXItem
TBXItem156Action)NonVisualDataModule.FullSynchronizeActionDisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem41  TTBXItem
TBXItem157Action!NonVisualDataModule.ConsoleAction  TTBXItem
TBXItem190ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem42  TTBXItem
TBXItem158Action.NonVisualDataModule.SynchronizeBrowsingAction2   TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem1Action)NonVisualDataModule.CheckForUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesActionOptions
tboDefault   TTBXSeparatorItemTBXSeparatorItem46  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft-Top� Caption   ÖverföringsinställningarDockPos,DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXLabelItemTransferSettingsLabelItemCaption   ÖverföringsinställningarMargin  TTBXDropDownItemTransferDropDown	EditWidth� Hint0   Välj förinställda överföringsinställningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelCaption    MarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarCustomCommandsToolbarLeft,Top� CaptionEgna kommandonChevronMenu	ChevronPriorityForNewItems
tbcpLowestDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrderVisible   �TPanelRemotePanelLeft�Top� Width�Height!Constraints.MinHeight� Constraints.MinWidth� ParentColor	TabOrder � 
TPathLabelRemotePathLabelLeft TopOWidth�HeightUnixPath	IndentVerticalAutoSizeVertical	HotTrack	OnGetStatusRemotePathLabelGetStatusOnPathClickRemotePathLabelPathClickOnMaskClickRemotePathLabelMaskClickAutoSizeTransparent
OnDblClickPathLabelDblClick  �	TSplitterRemotePanelSplitterLeft Top� Width�HeightCursorcrSizeNSHinti   Dra för att ändra storlek på katalogträd. Dubbelklicka för att gör höjden på katalogträden lika.AlignalTop  �TTBXStatusBarRemoteStatusBarTopWidth�PanelsFramedSize� StretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint    Klicka för att visa dolda filerMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint,   Klicka för att ändra eller ta bort filtretMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis  OnPanelClickRemoteStatusBarPanelClick  �TPanelRemoteDirPanelLeft Top� Width�HeightqConstraints.MinHeightF �TUnixDirViewRemoteDirViewWidthHeightq
NortonLikenlOnOnUpdateStatusBarRemoteDirViewUpdateStatusBar	PathLabelRemotePathLabelAddParentDir	OnDDFileOperationExecuted(RemoteFileControlDDFileOperationExecutedOnHistoryGoDirViewHistoryGoOnPathChangeRemoteDirViewPathChange  �TTBXToolbarReconnectToolbarTabOrder  TDirViewOtherLocalDirViewLeftTop Width� HeightqAlignalRightConstraints.MinHeightFDoubleBuffered	FullDrag	HideSelectionIconOptions.AutoArrange	ParentDoubleBuffered	PopupMenu&NonVisualDataModule.RemoteDirViewPopupTabOrderOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterOtherLocalDirViewEnterOnExitDirViewExit	OnKeyDownDirViewKeyDown
OnKeyPressDirViewKeyPressDirColProperties.ExtVisibleOnUpdateStatusBar OtherLocalDirViewUpdateStatusBarAddParentDir	OnSelectItemDirViewSelectItemOnLoadedDirViewLoadedOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDTargetHasDropHandler"LocalDirViewDDTargetHasDropHandlerOnDDFileOperationLocalFileControlDDFileOperation
OnExecFileLocalDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayDirViewGetOverlayConfirmDeleteUseIconUpdateThread	WatchForChanges	OnFileIconForNameLocalDirViewFileIconForNameOnContextPopupOtherLocalDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnHistoryGoDirViewHistoryGoOnPathChangeOtherLocalDirViewPathChangeOnBusyDirViewBusyOnChangeFocusDirViewChangeFocusDirViewStyle	dvsReport   �TPanelRemoteDrivePanelTopdWidth�Height-AlignalTopConstraints.MinHeight � 
TDriveViewOtherLocalDriveViewLeftTop Width� Height-WatchDirectory	DirViewOtherLocalDirViewOnRefreshDrivesLocalDriveViewRefreshDrivesOnBusyDirViewBusyOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDFileOperationLocalFileControlDDFileOperationAlignalRightConstraints.MinHeightDoubleBuffered	HideSelectionIndentParentColorParentDoubleBufferedTabOrderTabStopOnEnterOtherLocalDriveViewEnterOnNeedHiddenDirectories#LocalDriveViewNeedHiddenDirectories  �TUnixDriveViewRemoteDriveViewWidthHeight-TabStop   TTBXDockRemoteTopDockLeft Top Width�HeightOFixAlign	OnContextPopupDockContextPopup TTBXToolbarRemoteHistoryToolbarLeft TopCaption   FjärrhistorikDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemRemoteBackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemRemoteForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	   TTBXToolbarRemoteNavigationToolbarLeftPTopCaption   FjärrnavigeringDockPosHDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem165Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem
TBXItem166Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem
TBXItem167Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem
TBXItem168Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem37  TTBXItem
TBXItem132Action*NonVisualDataModule.RemoteFindFilesAction2DisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem44  TTBXItem
TBXItem170Action$NonVisualDataModule.RemoteTreeAction  TTBXSubmenuItemTBXSubmenuItem32Caption   Ändra stil för katalogvy
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem278Action&NonVisualDataModule.RemoteReportAction  TTBXSeparatorItemTBXSeparatorItem78  TTBXItem
TBXItem279Action)NonVisualDataModule.RemoteThumbnailAction    TTBXToolbarRemotePathToolbarLeft Top Caption   Fjärrsökväg
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemRemotePathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXSubmenuItemRemoteOpenDirButtonAction'NonVisualDataModule.RemoteOpenDirActionDropdownCombo	OnPopupRemoteOpenDirButtonPopup  TTBXSubmenuItem
TBXItem229Action&NonVisualDataModule.RemoteFilterActionDropdownCombo	 TTBXItem
TBXItem169Action&NonVisualDataModule.RemoteFilterActionOptions
tboDefault   TTBXSeparatorItemTBXSeparatorItem63  TTBXItem
TBXItem237Action/NonVisualDataModule.FileColorsPreferencesAction    TTBXToolbarRemoteFileToolbarLeftTop5Caption   FjärrfilerDockPosDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemRemoteCopyItemAction$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem143Action,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItem
TBXItem200Action)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem59  TTBXItemRemoteMoveItemAction$NonVisualDataModule.RemoteMoveAction   TTBXSeparatorItemTBXSeparatorItem55  TTBXSubmenuItem
TBXItem242Action%NonVisualDataModule.RemoteEditAction2DisplayModenbdmImageAndTextDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem
TBXItem241Action'NonVisualDataModule.RemoteDeleteAction2  TTBXItem
TBXItem240Action'NonVisualDataModule.RemoteRenameAction2  TTBXSubmenuItem
TBXItem243Action+NonVisualDataModule.RemotePropertiesAction2DisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem259Action+NonVisualDataModule.RemotePropertiesAction2Options
tboDefault   TTBXSeparatorItemTBXSeparatorItem71  TTBXItem
TBXItem260Action7NonVisualDataModule.RemoteCalculateDirectorySizesAction   TTBXSeparatorItemTBXSeparatorItem56  TTBXSubmenuItemRemoteNewSubmenuItemCaption&NyDisplayModenbdmImageAndTextHintSkapa objekt|Skapa nytt objekt
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem247Action'NonVisualDataModule.RemoteNewFileAction  TTBXItem
TBXItem244Action*NonVisualDataModule.RemoteCreateDirAction3  TTBXItem
TBXItem246Action,NonVisualDataModule.RemoteAddEditLinkAction3    TTBXToolbarRemoteSelectionToolbarLeftHTopCaption   FjärrmarkeringDockPosDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem138Action'NonVisualDataModule.RemoteSelectAction2  TTBXItem
TBXItem139Action)NonVisualDataModule.RemoteUnselectAction2  TTBXItem
TBXItem140Action*NonVisualDataModule.RemoteSelectAllAction2    TTBXDockRemoteBottomDockLeft TopWidth�Height	FixAlign	PositiondpBottom   �TPanel
QueuePanelTopWidth�HeighttParentColor	TabOrder �
TPathLabel
QueueLabelWidth�  �	TSplitterQueueFileListSplitterTop]Width�  �	TListView
QueueView3Width�Height.TabStop  �TTBXDock	QueueDockWidth�  �	TListViewQueueFileListTop`Width�   �TThemePageControlSessionsPageControlTop� Width�  �TPanel
LocalPanelLeft Top� Width�Height!AlignalLeft
BevelOuterbvNoneConstraints.MinHeight� Constraints.MinWidth� ParentBackgroundParentColor	TabOrder  
TPathLabelLocalPathLabelLeft TopOWidth�HeightIndentVerticalAutoSizeVertical	HotTrack	OnGetStatusLocalPathLabelGetStatusOnPathClickLocalPathLabelPathClickOnMaskClickLocalPathLabelMaskClickAutoSize	PopupMenu#NonVisualDataModule.LocalPanelPopupTransparent
OnDblClickPathLabelDblClick  	TSplitterLocalPanelSplitterLeft Top� Width�HeightCursorcrSizeNSHinti   Dra för att ändra storlek på katalogträd. Dubbelklicka för att gör höjden på katalogträden lika.AlignalTopAutoSnapMinSizeFResizeStylersUpdate  TTBXStatusBarLocalStatusBarLeft TopWidth�HeightPanelsFramedSize� StretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint    Klicka för att visa dolda filerMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaRightJustifyFramedHint,   Klicka för att ändra eller ta bort filtretMaxSizexSizePStretchPriorityTag TextTruncationtwEndEllipsis  ParentShowHintShowHint	UseSystemFontOnClickLocalStatusBarClickOnPanelClickLocalStatusBarPanelClick  TDirViewLocalDirViewLeft Top� Width�HeightqAlignalClientConstraints.MinHeightFDoubleBuffered	FullDrag	HideSelectionIconOptions.AutoArrange	ParentDoubleBuffered	PopupMenu%NonVisualDataModule.LocalDirViewPopupTabOrderOnColumnRightClickDirViewColumnRightClick	OnEditingDirViewEditingOnEnterLocalDirViewEnterOnExitDirViewExit	OnKeyDownDirViewKeyDown
OnKeyPressDirViewKeyPressDirColProperties.ExtVisible	PathLabelLocalPathLabelOnUpdateStatusBarLocalDirViewUpdateStatusBarAddParentDir	OnSelectItemDirViewSelectItemOnLoadedDirViewLoadedOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDTargetHasDropHandler"LocalDirViewDDTargetHasDropHandlerOnDDFileOperationLocalFileControlDDFileOperation
OnExecFileLocalDirViewExecFileOnMatchMaskDirViewMatchMaskOnGetOverlayDirViewGetOverlayConfirmDeleteUseIconUpdateThread	WatchForChanges	OnFileIconForNameLocalDirViewFileIconForNameOnContextPopupLocalDirViewContextPopupOnHistoryChangeDirViewHistoryChangeOnHistoryGoDirViewHistoryGoOnPathChangeLocalDirViewPathChangeOnBusyDirViewBusyOnChangeFocusDirViewChangeFocusDirViewStyle	dvsReport  TTBXDockLocalTopDockLeft Top Width�HeightOFixAlign	OnContextPopupDockContextPopup TTBXToolbarLocalHistoryToolbarLeft TopCaptionLokal historikDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemLocalBackButtonAction#NonVisualDataModule.LocalBackActionDropdownCombo	  TTBXSubmenuItemLocalForwardButtonAction&NonVisualDataModule.LocalForwardActionDropdownCombo	   TTBXToolbarLocalNavigationToolbarLeftPTopCaptionLokal navigeringDockPosDDockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem159Action(NonVisualDataModule.LocalParentDirAction  TTBXItem
TBXItem160Action&NonVisualDataModule.LocalRootDirAction  TTBXItem
TBXItem161Action&NonVisualDataModule.LocalHomeDirAction  TTBXItem
TBXItem162Action&NonVisualDataModule.LocalRefreshAction  TTBXSeparatorItemTBXSeparatorItem43  TTBXItem
TBXItem164Action#NonVisualDataModule.LocalTreeAction  TTBXSubmenuItemTBXSubmenuItem4Caption   Ändra stil för katalogvy
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem269Action%NonVisualDataModule.LocalReportAction  TTBXSeparatorItemTBXSeparatorItem75  TTBXItem
TBXItem268Action(NonVisualDataModule.LocalThumbnailAction    TTBXToolbarLocalPathToolbarLeft Top Caption   Lokal sökväg
DockableTodpTopdpBottom DockModedmCannotFloatDockPos ImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	Stretch	TabOrder OnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXComboBoxItemLocalPathComboBox	EditWidth� 	ShowImage	DropDownList	MaxVisibleItemsShowListImages	OnAdjustImageIndex!LocalPathComboBoxAdjustImageIndexOnItemClickLocalPathComboBoxItemClickOnCancelLocalPathComboBoxCancel  TTBXSubmenuItemLocalOpenDirButtonAction&NonVisualDataModule.LocalOpenDirActionDropdownCombo	OnPopupLocalOpenDirButtonPopup  TTBXSubmenuItem
TBXItem228Action%NonVisualDataModule.LocalFilterActionDropdownCombo	 TTBXItem
TBXItem245Action%NonVisualDataModule.LocalFilterAction  TTBXSeparatorItemTBXSeparatorItem64  TTBXItem
TBXItem251Action/NonVisualDataModule.FileColorsPreferencesAction    TTBXToolbarLocalFileToolbarLeft Top5CaptionLokala filerDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemLocalCopyItemAction#NonVisualDataModule.LocalCopyActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem144Action+NonVisualDataModule.LocalCopyNonQueueAction  TTBXItem
TBXItem174Action(NonVisualDataModule.LocalCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem58  TTBXItemLocalMoveItemAction#NonVisualDataModule.LocalMoveAction   TTBXSeparatorItemTBXSeparatorItem54  TTBXSubmenuItem
TBXItem235Action$NonVisualDataModule.LocalEditAction2DisplayModenbdmImageAndTextDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem
TBXItem234Action&NonVisualDataModule.LocalDeleteAction2  TTBXItem
TBXItem233Action&NonVisualDataModule.LocalRenameAction2  TTBXSubmenuItem
TBXItem236Action*NonVisualDataModule.LocalPropertiesAction2DisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem258Action*NonVisualDataModule.LocalPropertiesAction2Options
tboDefault   TTBXSeparatorItemTBXSeparatorItem70  TTBXItem
TBXItem113Action6NonVisualDataModule.LocalCalculateDirectorySizesAction   TTBXSeparatorItemTBXSeparatorItem35  TTBXSubmenuItemLocalNewSubmenuItemCaption&NyDisplayModenbdmImageAndTextHintSkapa objekt|Skapa nytt objekt
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem248Action&NonVisualDataModule.LocalNewFileAction  TTBXItem
TBXItem249Action)NonVisualDataModule.LocalCreateDirAction3  TTBXItem
TBXItem250Action+NonVisualDataModule.LocalAddEditLinkAction3    TTBXToolbarLocalSelectionToolbarLeft� TopCaptionLokal markeringDockPos� DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem137Action&NonVisualDataModule.LocalSelectAction2  TTBXItem	TBXItem32Action(NonVisualDataModule.LocalUnselectAction2  TTBXItem	TBXItem30Action)NonVisualDataModule.LocalSelectAllAction2    
TDriveViewLocalDriveViewLeft TopdWidth�Height-WatchDirectory	DirViewLocalDirViewOnRefreshDrivesLocalDriveViewRefreshDrivesOnBusyDirViewBusyOnDDDragEnterLocalFileControlDDDragEnterOnDDDragLeaveFileControlDDDragLeaveOnDDFileOperationLocalFileControlDDFileOperationAlignalTopConstraints.MinHeightDoubleBuffered	HideSelectionIndentParentColorParentDoubleBufferedTabOrderTabStopOnEnterLocalDriveViewEnterOnNeedHiddenDirectories#LocalDriveViewNeedHiddenDirectories  TTBXDockLocalBottomDockLeft TopWidth�Height	FixAlign	PositiondpBottom   �TTBXDock
BottomDockLeft Top�Width�Height5FixAlign	PositiondpBottomOnContextPopupDockContextPopup TTBXToolbarToolbar2ToolbarLeft TopCaptionSnabbtangenterDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHintStretch	TabOrder Visible TTBXItem
TBXItem171Action'NonVisualDataModule.CurrentRenameActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem172Action%NonVisualDataModule.CurrentEditActionDisplayModenbdmImageAndTextStretch	  TTBXItemCurrentCopyToolbar2ItemAction$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndTextStretch	  TTBXItemCurrentMoveToolbar2ItemAction$NonVisualDataModule.RemoteMoveActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem175Action*NonVisualDataModule.CurrentCreateDirActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem176Action'NonVisualDataModule.CurrentDeleteActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem177Action+NonVisualDataModule.CurrentPropertiesActionDisplayModenbdmImageAndTextStretch	  TTBXItem
TBXItem178Action+NonVisualDataModule.CloseApplicationAction2DisplayModenbdmImageAndTextStretch	   TTBXToolbarCommandLineToolbarLeft Top CaptionCommandLineToolbarDockModedmCannotFloatStretch	TabOrderVisibleOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize TTBXLabelItemCommandLinePromptLabelCaption
CommandX >Margin  TTBXComboBoxItemCommandLineComboOnBeginEditCommandLineComboBeginEditExtendedAccept	OnPopupCommandLineComboPopup    �TTBXStatusBar	StatusBarLeft Top�Width�ImagesGlyphsModule.SessionImagesPanelsSizedStretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  ParentShowHint	PopupMenu%NonVisualDataModule.CommanderBarPopupShowHint	UseSystemFontOnPanelDblClickStatusBarPanelDblClick  �	TPanelQueueSeparatorPanelLeft TopWidth�HeightAlignalBottom
BevelEdgesbeBottom 	BevelKindbkFlatTabOrder  �TTBXDockMessageDockTop� Width�  �TApplicationEventsApplicationEventsLeftHTop`     TPF0�TScpExplorerFormScpExplorerFormLeft� Top� HelpType	htKeywordHelpKeywordui_explorerActiveControlRemoteDirViewCaptionScpExplorerFormClientHeight�ClientWidthx
TextHeight �	TSplitterQueueSplitterTopLWidthx  �TTBXDockTopDockWidthxHeight� OnContextPopupDockContextPopup TTBXToolbarMenuToolbarLeft Top CaptionMenyCloseButtonImagesGlyphsModule.ExplorerImagesMenuBar	OptionstboNoAutoHinttboShowHint 
ShrinkModetbsmWrapStretch	TabOrder  TTBXSubmenuItemTBXSubmenuItem5Caption&FilHelpKeywordui_explorer_menu#filesHintFiloperationer TTBXSubmenuItemTBXSubmenuItem26Caption&NyHelpKeyword
task_indexHintSkapa objekt|Skapa nytt objekt TTBXItem
TBXItem135Action!NonVisualDataModule.NewFileAction  TTBXItem
TBXItem136Action NonVisualDataModule.NewDirAction  TTBXItem
TBXItem209Action!NonVisualDataModule.NewLinkAction   TTBXSeparatorItemTBXSeparatorItem20  TTBXItem	TBXItem25Action%NonVisualDataModule.CurrentOpenAction  TTBXSubmenuItem	TBXItem26Action%NonVisualDataModule.RemoteEditAction2DropdownCombo	OnPopupEditMenuItemPopup  TTBXItemTBXItem4Action,NonVisualDataModule.CurrentAddEditLinkAction  TTBXSeparatorItemTBXSeparatorItem7  TTBXItem	TBXItem34Action'NonVisualDataModule.RemoteDeleteAction2  TTBXItem	TBXItem35Action'NonVisualDataModule.RemoteRenameAction2  TTBXItem	TBXItem41Action+NonVisualDataModule.RemotePropertiesAction2  TTBXItem	TBXItem61Action1NonVisualDataModule.CalculateDirectorySizesAction  TTBXSeparatorItemTBXSeparatorItem8  TTBXSubmenuItem	TBXItem30Action$NonVisualDataModule.RemoteCopyActionDropdownCombo	 TTBXItem
TBXItem156Action,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItem
TBXItem158Action)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem39  TTBXItem	TBXItem32Action$NonVisualDataModule.RemoteMoveAction   TTBXItem	TBXItem31Action&NonVisualDataModule.RemoteCopyToAction  TTBXItem	TBXItem33Action&NonVisualDataModule.RemoteMoveToAction  TTBXSeparatorItemTBXSeparatorItem42  TTBXItem	TBXItem62Action1NonVisualDataModule.CurrentCopyToClipboardAction2  TTBXItem	TBXItem36Action NonVisualDataModule.PasteAction3  TTBXSeparatorItemTBXSeparatorItem9  TTBXSubmenuItemCustomCommandsMenuAction,NonVisualDataModule.CustomCommandsFileAction  TTBXSubmenuItemTBXSubmenuItem6Caption&FilnamnHelpKeyword	filenamesHint$   Operationer med namn på valda filer TTBXItem	TBXItem38Action-NonVisualDataModule.FileListToClipboardAction  TTBXItem	TBXItem39Action1NonVisualDataModule.FullFileListToClipboardAction  TTBXItem	TBXItem40Action*NonVisualDataModule.FileGenerateUrlAction2   TTBXSubmenuItemTBXSubmenuItem25Caption	   &LåsningHint   Hantera fillås TTBXItem
TBXItem214ActionNonVisualDataModule.LockAction  TTBXItem
TBXItem216Action NonVisualDataModule.UnlockAction   TTBXSeparatorItemTBXSeparatorItem1  TTBXItemTBXItem1Action"NonVisualDataModule.CloseTabAction  TTBXItemTBXItem2Action+NonVisualDataModule.CloseApplicationAction2   TTBXSubmenuItemTBXSubmenuItem7Caption
&KommandonHelpKeywordui_explorer_menu#commandsHintAndra kommandon TTBXItem	TBXItem43Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem44Action)NonVisualDataModule.FullSynchronizeAction  TTBXItemTBXItem3Action*NonVisualDataModule.RemoteFindFilesAction2  TTBXSubmenuItemQueueSubmenuItemCaption   &KöHelpKeywordui_queue#manageHint   Kommandon för kölistaOnPopupQueueSubmenuItemPopup TTBXItemQueueEnableItem2Action%NonVisualDataModule.QueueEnableAction  TTBXItem	TBXItem46Action#NonVisualDataModule.QueueGoToAction  TTBXSeparatorItemTBXSeparatorItem10  TTBXItem	TBXItem47Action(NonVisualDataModule.QueueItemQueryAction  TTBXItem	TBXItem48Action(NonVisualDataModule.QueueItemErrorAction  TTBXItem	TBXItem49Action)NonVisualDataModule.QueueItemPromptAction  TTBXSeparatorItemTBXSeparatorItem11  TTBXItem	TBXItem50Action*NonVisualDataModule.QueueItemExecuteAction  TTBXItem
TBXItem196Action(NonVisualDataModule.QueueItemPauseAction  TTBXItem
TBXItem197Action)NonVisualDataModule.QueueItemResumeAction  TTBXItem	TBXItem51Action)NonVisualDataModule.QueueItemDeleteAction  TTBXComboBoxItemQueueSpeedComboBoxItemAction(NonVisualDataModule.QueueItemSpeedAction  TTBXSeparatorItemTBXSeparatorItem12  TTBXItem	TBXItem52Action%NonVisualDataModule.QueueItemUpAction  TTBXItem	TBXItem53Action'NonVisualDataModule.QueueItemDownAction  TTBXSeparatorItemTBXSeparatorItem48  TTBXSubmenuItemTBXSubmenuItem13Caption&AllaHelpKeywordui_queue#manageHint&   Administrationskommandon för kömassa TTBXItem
TBXItem198Action'NonVisualDataModule.QueuePauseAllAction  TTBXItem
TBXItem199Action(NonVisualDataModule.QueueResumeAllAction  TTBXItem
TBXItem154Action(NonVisualDataModule.QueueDeleteAllAction  TTBXSeparatorItemTBXSeparatorItem35  TTBXItem
TBXItem143Action,NonVisualDataModule.QueueDeleteAllDoneAction    TTBXSubmenuItemTBXSubmenuItem28Action/NonVisualDataModule.CustomCommandsNonFileAction  TTBXSeparatorItemTBXSeparatorItem13  TTBXItemTBXItem5Action,NonVisualDataModule.RemoteAddBookmarkAction2  TTBXItemTBXItem6Action0NonVisualDataModule.RemotePathToClipboardAction2  TTBXSeparatorItemTBXSeparatorItem2  TTBXItem	TBXItem54Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem55ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem14  TTBXItem	TBXItem57Action%NonVisualDataModule.ClearCachesAction   TTBXSubmenuItemTBXSubmenuItem18Caption&MarkeraHelpKeywordui_explorer_menu#markHint   Kommandon för markera TTBXItem
TBXItem107Action#NonVisualDataModule.SelectOneAction  TTBXItem
TBXItem108Action NonVisualDataModule.SelectAction  TTBXItem
TBXItem109Action"NonVisualDataModule.UnselectAction  TTBXItem
TBXItem110Action#NonVisualDataModule.SelectAllAction  TTBXSeparatorItemTBXSeparatorItem41  TTBXItem
TBXItem111Action)NonVisualDataModule.InvertSelectionAction  TTBXItem
TBXItem112Action(NonVisualDataModule.ClearSelectionAction  TTBXItem	TBXItem27Action*NonVisualDataModule.RestoreSelectionAction  TTBXSeparatorItemTBXSeparatorItem61  TTBXItem
TBXItem212Action'NonVisualDataModule.SelectSameExtAction  TTBXItem
TBXItem213Action)NonVisualDataModule.UnselectSameExtAction   TTBXSubmenuItemTBXSubmenuItem29Caption&FlikarHelpKeywordui_explorer_menu#tabsHintFlikkommandon TTBXItem
TBXItem113Action NonVisualDataModule.NewTabAction  TTBXItem
TBXItem166Action"NonVisualDataModule.CloseTabAction  TTBXItem
TBXItem218Action&NonVisualDataModule.DuplicateTabAction  TTBXItem
TBXItem167Action#NonVisualDataModule.RenameTabAction  TTBXSeparatorItemTBXSeparatorItem47  TTBXColorItemColorMenuItemAction$NonVisualDataModule.ColorMenuAction2ColorclNone  TTBXSeparatorItemTBXSeparatorItem49  TTBXItem
TBXItem162Action+NonVisualDataModule.DisconnectSessionAction  TTBXItem
TBXItem163Action*NonVisualDataModule.ReconnectSessionAction  TTBXItem
TBXItem114Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem50  TTBXItem	TBXItem56Action(NonVisualDataModule.FileSystemInfoAction  TTBXItem
TBXItem144Action-NonVisualDataModule.SessionGenerateUrlAction2  TTBXItem
TBXItem160Action(NonVisualDataModule.ChangePasswordAction  TTBXItem	TBXItem14Action*NonVisualDataModule.PrivateKeyUploadAction  TTBXSeparatorItemTBXSeparatorItem37  TTBXSubmenuItemTBXSubmenuItem9Action$NonVisualDataModule.OpenedTabsAction  TTBXSubmenuItemTBXSubmenuItem10Action$NonVisualDataModule.WorkspacesAction  TTBXItem
TBXItem168Action'NonVisualDataModule.SaveWorkspaceAction  TTBXSeparatorItemTBXSeparatorItem53  TTBXSubmenuItemTBXSubmenuItem20Action(NonVisualDataModule.SavedSessionsAction2   TTBXSubmenuItemTBXSubmenuItem1Caption&VisaHelpKeywordui_explorer_menu#viewHint   Ändra layout för program TTBXSubmenuItemTBXSubmenuItem2Caption   &VerktygsfältHelpKeywordui_toolbarsHint   Visa/dölj verktygsfält TTBXItemTBXItem7Action-NonVisualDataModule.ExplorerAddressBandAction  TTBXItemTBXItem8Action-NonVisualDataModule.ExplorerToolbarBandAction  TTBXItemTBXItem9Action/NonVisualDataModule.ExplorerSelectionBandAction  TTBXItem	TBXItem10Action.NonVisualDataModule.ExplorerSessionBandAction2  TTBXItem	TBXItem11Action1NonVisualDataModule.ExplorerPreferencesBandAction  TTBXItem	TBXItem12Action*NonVisualDataModule.ExplorerSortBandAction  TTBXItem	TBXItem82Action-NonVisualDataModule.ExplorerUpdatesBandAction  TTBXItem	TBXItem83Action.NonVisualDataModule.ExplorerTransferBandAction  TTBXItem	TBXItem28Action4NonVisualDataModule.ExplorerCustomCommandsBandAction  TTBXSeparatorItemTBXSeparatorItem19  TTBXItem	TBXItem92Action&NonVisualDataModule.LockToolbarsAction  TTBXItem
TBXItem140Action.NonVisualDataModule.SelectiveToolbarTextAction  TTBXSubmenuItem
TBXItem169Action)NonVisualDataModule.ToolbarIconSizeAction TTBXItem
TBXItem273Action/NonVisualDataModule.ToolbarIconSizeNormalAction	RadioItem	  TTBXItem
TBXItem274Action.NonVisualDataModule.ToolbarIconSizeLargeAction	RadioItem	  TTBXItem
TBXItem275Action2NonVisualDataModule.ToolbarIconSizeVeryLargeAction	RadioItem	    TTBXItemSessionsTabs3Action'NonVisualDataModule.SessionsTabsAction2  TTBXItem	TBXItem13Action#NonVisualDataModule.StatusBarAction  TTBXSubmenuItemTBXSubmenuItem14Caption   &KöHelpKeywordui_queueHint   Konfigurera kölista TTBXItem	TBXItem77Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem	TBXItem78Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem	TBXItem79Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem21  TTBXItem	TBXItem80Action&NonVisualDataModule.QueueToolbarAction  TTBXItem
TBXItem164Action'NonVisualDataModule.QueueFileListAction  TTBXSeparatorItemTBXSeparatorItem51  TTBXItem
TBXItem115Action1NonVisualDataModule.QueueResetLayoutColumnsAction  TTBXSeparatorItemTBXSeparatorItem22  TTBXSubmenuItemTBXSubmenuItem8Action-NonVisualDataModule.QueueCycleOnceEmptyActionDropdownCombo	 TTBXItem
TBXItem222Action,NonVisualDataModule.QueueIdleOnceEmptyAction	RadioItem	  TTBXItem
TBXItem223Action3NonVisualDataModule.QueueDisconnectOnceEmptyAction2	RadioItem	  TTBXItem
TBXItem148Action0NonVisualDataModule.QueueSuspendOnceEmptyAction2  TTBXItem
TBXItem224Action1NonVisualDataModule.QueueShutDownOnceEmptyAction2	RadioItem	   TTBXItem	TBXItem81Action*NonVisualDataModule.QueuePreferencesAction   TTBXItem	TBXItem15Action$NonVisualDataModule.RemoteTreeAction  TTBXSeparatorItemTBXSeparatorItem3  TTBXItem	TBXItem16Action$NonVisualDataModule.RemoteIconAction  TTBXItem	TBXItem17Action)NonVisualDataModule.RemoteSmallIconAction  TTBXItem	TBXItem18Action$NonVisualDataModule.RemoteListAction  TTBXItem	TBXItem19Action&NonVisualDataModule.RemoteReportAction  TTBXItem
TBXItem170Action)NonVisualDataModule.RemoteThumbnailAction  TTBXSeparatorItemTBXSeparatorItem4  TTBXSubmenuItemTBXSubmenuItem15Caption	   &Gå tillHelpKeywordtask_navigateHint   Gå till katalog TTBXItem	TBXItem84Action'NonVisualDataModule.RemoteOpenDirAction  TTBXSeparatorItemTBXSeparatorItem25  TTBXItem	TBXItem85Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem86Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem87Action'NonVisualDataModule.RemoteHomeDirAction  TTBXSeparatorItemTBXSeparatorItem26  TTBXItem	TBXItem88Action$NonVisualDataModule.RemoteBackAction  TTBXItem	TBXItem89Action'NonVisualDataModule.RemoteForwardAction   TTBXItem	TBXItem20Action'NonVisualDataModule.RemoteRefreshAction  TTBXSubmenuItemTBXSubmenuItem16Caption&SorteraHelpKeywordui_file_panel#sorting_filesHint   Ändra filordning i panelen TTBXItem	TBXItem93Action.NonVisualDataModule.RemoteSortAscendingAction2  TTBXSeparatorItemTBXSeparatorItem28  TTBXItem	TBXItem94Action+NonVisualDataModule.RemoteSortByNameAction2
GroupIndex  TTBXItem	TBXItem95Action*NonVisualDataModule.RemoteSortByExtAction2
GroupIndex  TTBXItem	TBXItem97Action+NonVisualDataModule.RemoteSortBySizeAction2
GroupIndex  TTBXItem
TBXItem132Action+NonVisualDataModule.RemoteSortByTypeAction2	RadioItem	  TTBXItem	TBXItem96Action.NonVisualDataModule.RemoteSortByChangedAction2
GroupIndex  TTBXItem	TBXItem98Action-NonVisualDataModule.RemoteSortByRightsAction2
GroupIndex  TTBXItem	TBXItem99Action,NonVisualDataModule.RemoteSortByOwnerAction2
GroupIndex  TTBXItem
TBXItem100Action,NonVisualDataModule.RemoteSortByGroupAction2
GroupIndex   TTBXSubmenuItemColumndsSubmenuItemCaption	&KolumnerHelpKeywordui_file_panel#selecting_columns TTBXItem
TBXItem101Action3NonVisualDataModule.ShowHideRemoteNameColumnAction2  TTBXItem
TBXItem102Action3NonVisualDataModule.ShowHideRemoteSizeColumnAction2  TTBXItem
TBXItem131Action3NonVisualDataModule.ShowHideRemoteTypeColumnAction2  TTBXItem
TBXItem103Action6NonVisualDataModule.ShowHideRemoteChangedColumnAction2  TTBXItem
TBXItem104Action5NonVisualDataModule.ShowHideRemoteRightsColumnAction2  TTBXItem
TBXItem105Action4NonVisualDataModule.ShowHideRemoteOwnerColumnAction2  TTBXItem
TBXItem106Action4NonVisualDataModule.ShowHideRemoteGroupColumnAction2  TTBXItem	TBXItem76Action9NonVisualDataModule.ShowHideRemoteLinkTargetColumnAction2  TTBXSeparatorItemTBXSeparatorItem73  TTBXItem
TBXItem264Action/NonVisualDataModule.AutoSizeRemoteColumnsAction  TTBXItem
TBXItem266Action2NonVisualDataModule.ResetLayoutRemoteColumnsAction   TTBXItem
TBXItem138Action&NonVisualDataModule.RemoteFilterAction  TTBXSeparatorItemTBXSeparatorItem5  TTBXItem	TBXItem21Action%NonVisualDataModule.PreferencesAction   TTBXSubmenuItemTBXSubmenuItem22Caption   &HjälpHelpKeywordui_explorer_menu#helpHint   Hjälp TTBXItem
TBXItem116Action)NonVisualDataModule.TableOfContentsAction  TTBXItem
TBXItem159ActionNonVisualDataModule.TipsAction  TTBXSeparatorItemTBXSeparatorItem30  TTBXItem
TBXItem117Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem118Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem119Action%NonVisualDataModule.HistoryPageAction  TTBXSeparatorItemTBXSeparatorItem31  TTBXItem
TBXItem120Action)NonVisualDataModule.CheckForUpdatesAction  TTBXSeparatorItemTBXSeparatorItem32  TTBXItem
TBXItem121Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem33  TTBXItem
TBXItem122ActionNonVisualDataModule.AboutAction    TTBXToolbarButtonsToolbarLeft Top4Caption	KommandonDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItem
BackButtonAction$NonVisualDataModule.RemoteBackActionDropdownCombo	  TTBXSubmenuItemForwardButtonAction'NonVisualDataModule.RemoteForwardActionDropdownCombo	  TTBXSeparatorItemTBXSeparatorItem6  TTBXItem	TBXItem23Action)NonVisualDataModule.RemoteParentDirAction  TTBXItem	TBXItem24Action'NonVisualDataModule.RemoteRootDirAction  TTBXItem	TBXItem29Action'NonVisualDataModule.RemoteHomeDirAction  TTBXItem	TBXItem37Action'NonVisualDataModule.RemoteRefreshAction  TTBXSeparatorItemTBXSeparatorItem24  TTBXItem
TBXItem139Action*NonVisualDataModule.RemoteFindFilesAction2DisplayModenbdmImageAndText  TTBXSeparatorItemTBXSeparatorItem15  TTBXSubmenuItem
TBXItem141Action$NonVisualDataModule.RemoteCopyActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem155Action,NonVisualDataModule.RemoteCopyNonQueueAction  TTBXItem
TBXItem157Action)NonVisualDataModule.RemoteCopyQueueAction  TTBXSeparatorItemTBXSeparatorItem38  TTBXItem
TBXItem142Action$NonVisualDataModule.RemoteMoveAction   TTBXSeparatorItemTBXSeparatorItem27  TTBXSubmenuItem	TBXItem42Action%NonVisualDataModule.RemoteEditAction2DisplayModenbdmImageAndTextDropdownCombo	OnPopupEditMenuItemPopup  TTBXItem	TBXItem45Action%NonVisualDataModule.CurrentOpenAction  TTBXItem	TBXItem58Action'NonVisualDataModule.RemoteDeleteAction2  TTBXSubmenuItem	TBXItem59Action+NonVisualDataModule.RemotePropertiesAction2DisplayModenbdmImageAndTextDropdownCombo	 TTBXItem	TBXItem90Action+NonVisualDataModule.RemotePropertiesAction2Options
tboDefault   TTBXSeparatorItemTBXSeparatorItem29  TTBXItem	TBXItem22Action7NonVisualDataModule.RemoteCalculateDirectorySizesAction   TTBXItem	TBXItem60Action'NonVisualDataModule.RemoteRenameAction2  TTBXSeparatorItemTBXSeparatorItem16  TTBXSubmenuItemNewSubmenuItemCaption&NyDisplayModenbdmImageAndTextHintSkapa objekt|Skapa nytt objekt
ImageIndexOptionstboDropdownArrow  TTBXItem
TBXItem247Action'NonVisualDataModule.RemoteNewFileAction  TTBXItem
TBXItem244Action*NonVisualDataModule.RemoteCreateDirAction3  TTBXItem
TBXItem246Action,NonVisualDataModule.RemoteAddEditLinkAction3   TTBXItem	TBXItem63Action!NonVisualDataModule.ConsoleAction  TTBXItem	TBXItem91ActionNonVisualDataModule.PuttyAction  TTBXSeparatorItemTBXSeparatorItem17  TTBXItem	TBXItem64Action%NonVisualDataModule.SynchronizeAction  TTBXItem	TBXItem65Action)NonVisualDataModule.FullSynchronizeActionDisplayModenbdmImageAndText   TTBXToolbarSelectionToolbarLeft TopNCaption	MarkeringDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem	TBXItem66Action NonVisualDataModule.SelectAction  TTBXItem	TBXItem67Action"NonVisualDataModule.UnselectAction  TTBXSeparatorItemTBXSeparatorItem18  TTBXItem	TBXItem68Action#NonVisualDataModule.SelectAllAction  TTBXItem	TBXItem69Action)NonVisualDataModule.InvertSelectionAction  TTBXItem	TBXItem70Action(NonVisualDataModule.ClearSelectionAction  TTBXItem
TBXItem134Action*NonVisualDataModule.RestoreSelectionAction   TTBXToolbarSessionToolbar2Left TophCaptionSessioner och flikarDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem123Action NonVisualDataModule.NewTabActionDisplayModenbdmImageAndText  TTBXItem
TBXItem125Action-NonVisualDataModule.SaveCurrentSessionAction2  TTBXSeparatorItemTBXSeparatorItem23  TTBXItem
TBXItem137Action&NonVisualDataModule.DuplicateTabAction  TTBXItem
TBXItem124Action"NonVisualDataModule.CloseTabAction  TTBXSeparatorItemTBXSeparatorItem34  TTBXSubmenuItemTBXSubmenuItem23Action(NonVisualDataModule.SavedSessionsAction2DisplayModenbdmImageAndTextOptionstboDropdownArrow    TTBXToolbarPreferencesToolbarLeft Top� Caption   InställningarDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem126Action%NonVisualDataModule.PreferencesAction  TTBXSeparatorItemTBXSeparatorItem36  TTBXSubmenuItemTBXSubmenuItem3Action*NonVisualDataModule.RemoteCycleStyleActionDropdownCombo	 TTBXItem	TBXItem72Action$NonVisualDataModule.RemoteIconAction  TTBXItem	TBXItem73Action)NonVisualDataModule.RemoteSmallIconAction  TTBXItem	TBXItem74Action$NonVisualDataModule.RemoteListAction  TTBXItem	TBXItem75Action&NonVisualDataModule.RemoteReportAction  TTBXItem
TBXItem279Action)NonVisualDataModule.RemoteThumbnailAction   TTBXSubmenuItemTBXSubmenuItem24Action)NonVisualDataModule.QueueToggleShowActionDisplayModenbdmImageAndTextDropdownCombo	 TTBXItem
TBXItem128Action#NonVisualDataModule.QueueShowAction	RadioItem	  TTBXItem
TBXItem129Action,NonVisualDataModule.QueueHideWhenEmptyAction	RadioItem	  TTBXItem
TBXItem130Action#NonVisualDataModule.QueueHideAction	RadioItem	  TTBXSeparatorItemTBXSeparatorItem44  TTBXItem
TBXItem165Action'NonVisualDataModule.QueueFileListAction   TTBXItem	TBXItem71Action$NonVisualDataModule.RemoteTreeAction   TTBXToolbarSortToolbarLeft Top� CaptionSorteraDockPos DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXItem
TBXItem145Action.NonVisualDataModule.CurrentSortAscendingAction  TTBXSeparatorItemTBXSeparatorItem40  TTBXItem
TBXItem146Action+NonVisualDataModule.CurrentSortByNameAction  TTBXItem
TBXItem147Action*NonVisualDataModule.CurrentSortByExtAction  TTBXItem
TBXItem133Action,NonVisualDataModule.CurrentSortByTypeAction2  TTBXItem
TBXItem149Action.NonVisualDataModule.CurrentSortByChangedAction  TTBXItem
TBXItem150Action+NonVisualDataModule.CurrentSortBySizeAction  TTBXItem
TBXItem151Action-NonVisualDataModule.CurrentSortByRightsAction  TTBXItem
TBXItem152Action,NonVisualDataModule.CurrentSortByOwnerAction  TTBXItem
TBXItem153Action,NonVisualDataModule.CurrentSortByGroupAction   TTBXToolbarAddressToolbarLeft TopCaptionAdress
DockableTodpTopdpBottom DockModedmCannotFloatDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHint	PopupMenu&NonVisualDataModule.RemoteAddressPopup	ResizableShowHint	Stretch	TabOrderOnResizeToolBarResizeOnGetBaseSizeToolbarGetBaseSize
OnEndModalAddressToolbarEndModal TTBXLabelItemTBXLabelItem1CaptionAdressMargin  TTBXComboBoxItemUnixPathComboBox	EditWidth� OnAcceptTextUnixPathComboBoxAcceptTextOnBeginEditUnixPathComboBoxBeginEdit	ShowImage	MaxVisibleItemsShowListImages	OnAdjustImageIndex"RemotePathComboBoxAdjustImageIndex
OnDrawItemRemotePathComboBoxDrawItemOnItemClickRemotePathComboBoxItemClickOnMeasureWidthRemotePathComboBoxMeasureWidthOnCancelRemotePathComboBoxCancel  TTBXSubmenuItemRemoteOpenDirButtonAction'NonVisualDataModule.RemoteOpenDirActionDropdownCombo	OnPopupRemoteOpenDirButtonPopup  TTBXSubmenuItem
TBXItem229Action&NonVisualDataModule.RemoteFilterActionDropdownCombo	 TTBXItem
TBXItem127Action&NonVisualDataModule.RemoteFilterAction  TTBXSeparatorItemTBXSeparatorItem43  TTBXItem
TBXItem161Action/NonVisualDataModule.FileColorsPreferencesAction    TTBXToolbarUpdatesToolbarLeft Top� CaptionUppdateringarDockPos�DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXSubmenuItemTBXSubmenuItem4Action)NonVisualDataModule.CheckForUpdatesActionDropdownCombo	 TTBXItem
TBXItem184Action)NonVisualDataModule.CheckForUpdatesActionOptions
tboDefault   TTBXSeparatorItemTBXSeparatorItem46  TTBXItem
TBXItem180Action"NonVisualDataModule.HomepageAction  TTBXItem
TBXItem187Action&NonVisualDataModule.DownloadPageAction  TTBXItem
TBXItem181Action#NonVisualDataModule.ForumPageAction  TTBXItem
TBXItem182Action%NonVisualDataModule.HistoryPageAction  TTBXItem
TBXItem185Action$NonVisualDataModule.DonatePageAction  TTBXSeparatorItemTBXSeparatorItem45  TTBXItem
TBXItem183Action,NonVisualDataModule.UpdatesPreferencesAction    TTBXToolbarTransferToolbarLeft-Top� Caption   ÖverföringsinställningarDockPos,DockRowImagesGlyphsModule.ExplorerImagesOptionstboShowHint ParentShowHintShowHint	TabOrder TTBXLabelItemTransferSettingsLabelItemCaption   ÖverföringsinställningarMargin  TTBXDropDownItemTransferDropDown	EditWidth� Hint0   Välj förinställda överföringsinställningarDropDownList	 TTBXStringListTransferListMaxVisibleItemsMinWidth^  TTBXLabelItemTransferLabelCaption    MarginShowAccelChar  TTBXSeparatorItemTBXSeparatorItem52  TTBXItem
TBXItem189Action,NonVisualDataModule.PresetsPreferencesActionDisplayModenbdmImageAndText    TTBXToolbarCustomCommandsToolbarLeft,Top� CaptionEgna kommandonChevronMenu	ChevronPriorityForNewItems
tbcpLowestDockPos� DockRowImagesGlyphsModule.ExplorerImagesParentShowHintShowHint	TabOrder	Visible   �TPanelRemotePanelLeft	Top� WidthfHeight]Constraints.MinHeight\Constraints.MinWidth�  �	TSplitterRemotePanelSplitterHeight>HintW   Dra för att ändra storlek på katalogträd. Dubbelklicka för att dölja katalogträd  �TTBXStatusBarRemoteStatusBarTopGWidthfHeightImagesGlyphsModule.SessionImagesPanelsSize� StretchPriorityTag TextTruncationtwEndEllipsis 	AlignmenttaCenterHint    Klicka för att visa dolda filerSizexTag TextTruncationtwEndEllipsis 	AlignmenttaCenterHint,   Klicka för att ändra eller ta bort filtretSizexTag TextTruncationtwEndEllipsis 	AlignmenttaCenterMaxSizeFViewPrioritybSizeFTag TextTruncationtwEndEllipsis 	AlignmenttaCenter
ImageIndexMaxSize#Size#Tag  	AlignmenttaCenterMaxSizePViewPrioritycSizePTag TextTruncationtwEndEllipsis  OnPanelClickRemoteStatusBarPanelClickOnPanelDblClickStatusBarPanelDblClick  �TPanelRemoteDirPanelWidth�Height> �TUnixDirViewRemoteDirViewWidth�Height>OnUpdateStatusBarRemoteDirViewUpdateStatusBarOnPathChangeRemoteDirViewPathChange   �TPanelRemoteDrivePanelHeight>Constraints.MinWidth( �TUnixDriveViewRemoteDriveViewHeight>   TTBXDock
BottomDockLeft Top>WidthfHeight	Color	clBtnFaceFixAlign	PositiondpBottom   �TPanel
QueuePanelTopOWidthx �
TPathLabel
QueueLabelWidthx  �	TSplitterQueueFileListSplitterWidthx  �	TListView
QueueView3Widthx  �TTBXDock	QueueDockWidthx  �	TListViewQueueFileListWidthx   �TThemePageControlSessionsPageControlTop� Widthx  �TTBXDockLeftDockLeft Top� Width	Height]PositiondpLeft  �TTBXDock	RightDockLeftoTop� Width	Height]PositiondpRight  �TTBXDockMessageDockTop� Widthx   TPF0TSelectMaskDialogSelectMaskDialogLeftqTopHelpType	htKeywordHelpKeyword	ui_selectBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSelectXClientHeight� ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style Position
poDesignedOnCloseQueryFormCloseQueryOnShowFormShow
DesignSize��  
TextHeight 	TGroupBox	MaskGroupLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize��   TLabelLabel3Left	Top	Width4HeightCaption	Fil&mask:FocusControlMaskEdit  TLabelColorFileNamesLabelLeft	TopMWidth� Height/AnchorsakLeftakTopakBottom AutoSizeCaption!about.html
index.html
photo.jpgColorclWindowParentColorShowAccelCharTransparentWordWrap	  TLabelColorSizesLabelLeft� TopMWidthRHeight/	AlignmenttaRightJustifyAnchorsakLeftakTopakBottom AutoSizeCaptionColorSizesLabelColorclWindowParentColorShowAccelCharTransparentWordWrap	  TLabelColorPaddingLabelLeft TopMWidth^Height/	AlignmenttaRightJustifyAnchorsakLeftakTopakRightakBottom AutoSizeColorclWindowParentColorShowAccelCharTransparentWordWrap	  	TCheckBoxApplyToDirectoriesCheckLeftTop6Width� HeightCaption   Tillämpa på &katalogerTabOrder  THistoryComboBoxMaskEditLeft	TopWidthUHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder Text*.*OnChangeMaskEditChangeOnExitMaskEditExit  TStaticTextHintTextLeft� Top0WidthsHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption	Mask&tipsTabOrderTabStop	  TButton
MaskButtonLeftdTopWidthPHeightAnchorsakTopakRight Caption	&RedigeraTabOrderOnClickMaskButtonClick  TButtonColorButtonLeftdTopMWidthPHeightAnchorsakTopakRight Caption   &FärgTabOrderOnClickColorButtonClick   TButtonOKBtnLeft� Top� WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeftTop� WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLefttTop� WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonClearButtonLeftrTop� WidthPHeightAnchorsakRightakBottom Caption&RensaModalResultTabOrderOnClickClearButtonClick   TPF0TSiteAdvancedDialogSiteAdvancedDialogLeft_Top� HelpType	htKeywordHelpKeywordui_login_advancedBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption"   Avancerade webbplatsinställningarClientHeight�ClientWidthkColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnClose	FormCloseOnCloseQueryFormCloseQueryOnShowFormShow
DesignSizek� 
TextHeight TPanel	MainPanelLeft Top WidthkHeight�AlignalTopAnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  TPageControlPageControlLeft� Top Width�Height�HelpType	htKeyword
ActivePageEnvironmentSheetAlignalClient	MultiLine	Style	tsButtonsTabOrderTabStopOnChangePageControlChange 	TTabSheetEnvironmentSheetTagHelpType	htKeywordHelpKeywordui_login_environmentCaption   Miljö
ImageIndex
TabVisible
DesignSize��  	TGroupBoxEnvironmentGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   ServermiljöTabOrder 
DesignSize��   TLabelEOLTypeLabelLeft	TopWidthHeightCaption1   Slut på rad &tecken (om det inte ges av server):FocusControlEOLTypeCombo  TLabelUtfLabelLeft	Top3Width� HeightCaption   &UTF-8 kodning på filnamn:FocusControlUtfCombo  TLabelTimeDifferenceLabelLeft	TopPWidth[HeightCaptionOffset tidszon:FocusControlTimeDifferenceEdit  TLabelTimeDifferenceHoursLabelLeft� TopPWidthHeightAnchorsakTopakRight CaptiontimmarFocusControlTimeDifferenceEdit  TLabelTimeDifferenceMinutesLabelLeftxTopPWidth+HeightAnchorsakTopakRight CaptionminuterFocusControlTimeDifferenceMinutesEdit  	TComboBoxEOLTypeComboLeftjTopWidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrder Items.StringsLFCR/LF   	TComboBoxUtfComboLeftjTop0WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrder  TUpDownEditTimeDifferenceEditLeft� TopMWidthLHeight	AlignmenttaRightJustifyMaxValue       �@MinValue       ��Value       ��AnchorsakTopakRight TabOrderOnChange
DataChange  TUpDownEditTimeDifferenceMinutesEditLeft&TopMWidthLHeight	AlignmenttaRightJustify	Increment       �@MaxValue       �@MinValue       ��Value       ��AnchorsakTopakRight TabOrderOnChange
DataChange  	TCheckBoxTimeDifferenceAutoCheckLeft� TopjWidthHeightAnchorsakTopakRight CaptionIdentifiera &automatisktTabOrderOnClick
DataChange  	TCheckBoxTrimVMSVersionsCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight CaptionTrimma VMS-versionsnummerTabOrderOnClick
DataChange   	TGroupBoxDSTModeGroupLeftTop� Width�Height]AnchorsakLeftakTopakRight Caption	SommartidTabOrder
DesignSize�]  TRadioButtonDSTModeUnixCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption7   Justera fjärrtidsstämpel med lokal ko&nvention (Unix)TabOrder OnClick
DataChange  TRadioButtonDSTModeWinCheckLeftTop.Width�HeightAnchorsakLeftakTopakRight Caption-   Justera fjärrtidsstämpel med &DST (Windows)TabOrderOnClick
DataChange  TRadioButtonDSTModeKeepCheckLeftTopEWidth�HeightAnchorsakLeftakTopakRight Caption    Bevara fjärrtidsstämpel (Unix)TabOrderOnClick
DataChange   	TGroupBox
PuttyGroupLeftTopWidth�HeightgAnchorsakLeftakTopakRight CaptionPuTTYTabOrder
DesignSize�g  TLabelPuttySettingsLabelLeft	TopWidth� HeightCaption   &PuTTY terminalinställningar:FocusControlEncryptKeyPasswordEdit  TButtonPuttySettingsButtonLeft	TopEWidth� HeightAnchorsakTopakRight Caption&Redigera i PuTTY...TabOrderOnClickPuttySettingsButtonClick  TEditPuttySettingsEditLeft	Top(Width�HeightAnchorsakLeftakTopakRight 	MaxLength@TabOrder TextPuttySettingsEditOnChange
DataChangeOnExitEncryptKeyEditExit    	TTabSheetDirectoriesSheetTagHelpType	htKeywordHelpKeywordui_login_directoriesCaption	Kataloger
ImageIndex
TabVisible
DesignSize��  	TGroupBoxDirectoriesGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize��   TLabelLocalDirectoryLabelLeft	TopsWidthQHeightCaption&Lokal katalogFocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft	TopDWidth^HeightCaption   F&järrkatalogFocusControlRemoteDirectoryEdit  TLabelLocalDirectoryDescLabelLeft	Top� WidthHeightCaptionB   Lokal katalog används inte i det utforskar-liknande gränssnittetShowAccelChar  TDirectoryEditLocalDirectoryEditLeft	Top� Width�HeightAcceptFiles	
DialogText    Välj lokal katalog vid uppstartClickKey@AnchorsakLeftakTopakRight TabOrderTextLocalDirectoryEditOnChange
DataChange  TEditRemoteDirectoryEditLeft	TopVWidth�HeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChange
DataChange  	TCheckBoxUpdateDirectoriesCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption"   Ko&m ihåg senast använda katalogTabOrder  	TCheckBoxSynchronizeBrowsingCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Syn&kronisera bläddringTabOrder    	TGroupBoxDirectoryOptionsGroupLeftTop� Width�HeighttAnchorsakLeftakTopakRight Caption   Alternativ vid kalalogläsningTabOrder
DesignSize�t  	TCheckBoxCacheDirectoriesCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Cacha &besökta fjärrkatalogerTabOrder OnClick
DataChange  	TCheckBoxCacheDirectoryChangesCheckLeftTop-WidthHeightAnchorsakLeftakTopakRight Caption   Cacha katalogf&örändringarTabOrderOnClick
DataChange  	TCheckBoxResolveSymlinksCheckLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption   Slå upp symboliska lä&nkarTabOrder  	TCheckBoxPreserveDirectoryChangesCheckLeft
Top-Width� HeightAnchorsakTopakRight Caption&Permanent cacheTabOrder  	TCheckBoxFollowDirectorySymlinksCheckLeftTop[Width�HeightAnchorsakLeftakTopakRight Caption(   &Följ symboliska länkar till katalogerTabOrder    	TTabSheetRecycleBinSheetTagHelpType	htKeywordHelpKeywordui_login_recycle_binCaptionPapperskorg
ImageIndex
TabVisible
DesignSize��  	TGroupBoxRecycleBinGroupLeftTopWidth�HeightwAnchorsakLeftakTopakRight CaptionPapperskorgTabOrder 
DesignSize�w  TLabelRecycleBinPathLabelLeft	TopDWidthhHeightCaption   Papp&erskorg på servernFocusControlRecycleBinPathEdit  	TCheckBoxDeleteToRecycleBinCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption6   Flytta borttagna filer på servern till &papperskorgenTabOrder OnClick
DataChange  	TCheckBoxOverwrittenToRecycleBinCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight CaptionG   Flytta &överskrivna filer på servern till papperskorgen (endast SFTP)TabOrderOnClick
DataChange  TEditRecycleBinPathEditLeft	TopVWidth�HeightAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRecycleBinPathEditOnChange
DataChange    	TTabSheetEncryptionSheetTagHelpType	htKeywordHelpKeywordui_login_encryptionCaption
Kryptering
TabVisible
DesignSize��  	TCheckBoxEncryptFilesCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption&Kryptera filerTabOrder OnClick
DataChange  	TGroupBoxEncryptFilesGroupLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   KrypteringsinställningarTabOrder
DesignSize�  TLabelLabel13Left	TopWidthQHeightCaptionKrypterings&nyckelFocusControlEncryptKeyPasswordEdit  TEditEncryptKeyVisibleEditLeft	Top(Width�HeightAnchorsakLeftakTopakRight 	MaxLength@TabOrderTextEncryptKeyVisibleEditVisibleOnChange
DataChangeOnExitEncryptKeyEditExit  TPasswordEditEncryptKeyPasswordEditLeft	Top(Width�HeightAnchorsakLeftakTopakRight 	MaxLength@TabOrder TextEncryptKeyPasswordEditOnChange
DataChangeOnExitEncryptKeyEditExit  	TCheckBoxShowEncryptionKeyCheckLeftTopEWidth�HeightCaption&Visa nyckelTabOrderOnClickShowEncryptionKeyCheckClick  TButtonGenerateKeyButtonLeft	Top\Width� HeightCaption&Generera nyckelTabOrderOnClickGenerateKeyButtonClick    	TTabSheet	SftpSheetTagHelpType	htKeywordHelpKeywordui_login_sftpCaptionSFTP
ImageIndex
TabVisible
DesignSize��  	TGroupBoxSFTPBugsGroupBoxLeftTop� Width�HeightMAnchorsakLeftakTopakRight Caption    Upptäckta buggar i SFTP servrarTabOrder
DesignSize�M  TLabelLabel10Left	TopWidth� HeightCaption;   &Omvänd ordning på symboliska länkar i kommandoargument:FocusControlSFTPBugSymlinkCombo  TLabelLabel36Left	Top/Width� HeightCaption3   Feltolkning av filtidsstä&mplar tidigare än 1970:FocusControlSFTPBugSignedTSCombo  	TComboBoxSFTPBugSymlinkComboLeftjTopWidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TComboBoxSFTPBugSignedTSComboLeftjTop,WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrder   	TGroupBoxSFTPProtocolGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize��   TLabelLabel34Left	Top3Width� HeightCaption"   Före&drar SFTP protokoll version:FocusControlSFTPMaxVersionCombo  TLabelLabel23Left	TopWidth?HeightCaptionSFTP ser&verFocusControlSftpServerEdit  TLabelLabel5Left	TopPWidth� HeightCaption"   &Kanonisera sökvägar på servernFocusControlSFTPRealPathCombo  	TComboBoxSFTPMaxVersionComboLeftjTop0WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderItems.StringsAuto0123456   	TComboBoxSftpServerEditLeft� TopWidthHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextSftpServerEditOnChange
DataChangeItems.StringsStandard/bin/sftp-serversudo su -c /bin/sftp-server   	TCheckBoxAllowScpFallbackCheckLeftTopjWidth�HeightAnchorsakLeftakTopakRight Caption   Tillåt SCP &fallbackTabOrderOnClick
DataChange  	TComboBoxSFTPRealPathComboLeftjTopMWidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrder  	TCheckBoxUsePosixRenameCheckLeftTop� Width�HeightAnchorsakLeftakTopakRight Caption   &Använd POSIX renameTabOrderOnClick
DataChange    	TTabSheetScpSheetTagHelpType	htKeywordHelpKeywordui_login_scpCaption
SCP/ShellX
ImageIndex
TabVisible
DesignSize��  	TGroupBoxOtherShellOptionsGroupLeftTop� Width�HeightHAnchorsakLeftakTopakRight Caption   Övriga alternativTabOrder
DesignSize�H  	TCheckBoxLookupUserGroupsCheckLeftTopWidth� HeightAllowGrayed	Caption   Slå upp &användargrupperTabOrder OnClick
DataChange  	TCheckBoxClearAliasesCheckLeftTop-Width� HeightCaptionRensa a&liasTabOrderOnClick
DataChange  	TCheckBoxUnsetNationalVarsCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight CaptionRensa &nationella variablerTabOrderOnClick
DataChange  	TCheckBoxScp1CompatibilityCheckLeft� Top-Width� HeightAnchorsakLeftakTopakRight Caption%   Använd scp&2 med scp1 kompatibilitetTabOrderOnClick
DataChange   	TGroupBox
ShellGroupLeftTopWidth�HeightQAnchorsakLeftakTopakRight CaptionSkalTabOrder 
DesignSize�Q  TLabelLabel19Left	TopWidthHeightCaptionS&kal:FocusControl	ShellEdit  TLabelLabel20Left	Top3WidthoHeightCaption&Returnera kodvariabel:FocusControlReturnVarEdit  	TComboBox	ShellEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrder Text	ShellEditItems.StringsStandard	/bin/bash/bin/ksh/bin/sh	sudo su -   	TComboBoxReturnVarEditLeft� Top0Width� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrderTextReturnVarEditItems.StringsAutomatisk identifiering?status    	TGroupBoxScpLsOptionsGroupLeftTopYWidth�HeightKAnchorsakLeftakTopakRight CaptionListning av katalogerTabOrder
DesignSize�K  TLabelLabel9Left	TopWidth`HeightCaption   &Kommando för listning:FocusControlListingCommandEdit  	TCheckBoxIgnoreLsWarningsCheckLeftTop0Width� HeightCaptionIgnorera LS &varningarTabOrderOnClick
DataChange  	TCheckBoxSCPLsFullTimeAutoCheckLeft� Top0Width� HeightAnchorsakLeftakTopakRight Caption#   Försök att få &full tidsstämpelTabOrderOnClick
DataChange  	TComboBoxListingCommandEditLeft� TopWidth� HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength2TabOrder TextListingCommandEditItems.Stringsls -lals -gla     	TTabSheetFtpSheetTagHelpType	htKeywordHelpKeywordui_login_ftpCaptionFTP
ImageIndex
TabVisible
DesignSize��  	TGroupBoxFtpGroupLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�  TLabelLabel25Left	Top0WidthwHeightCaption&Kommandon efter inloggning:FocusControlPostLoginCommandsMemo  TLabelFtpListAllLabelLeft	Top� Width� HeightCaption%   &Support för listning av dolda filerFocusControlFtpListAllCombo  TLabelLabel24Left	Top� Width� HeightCaption,   Använd &MLSD kommandon för kataloglistningFocusControlFtpUseMlsdCombo  TLabelFtpForcePasvIpLabelLeft	Top� Width� HeightCaption+   &Tvinga ip-adress för passiva anslutningarFocusControlFtpForcePasvIpCombo  TLabelFtpAccountLabelLeft	TopWidth0HeightCaptionK&onto:FocusControlFtpAccountEdit  TLabelLabel3Left	Top� Width� HeightCaption8   Använd &HOST-kommando för att välja värd på servernFocusControlFtpHostCombo  TMemoPostLoginCommandsMemoLeft	TopBWidth�Height5AnchorsakLeftakTopakRight 
ScrollBars
ssVerticalTabOrder  	TComboBoxFtpListAllComboLeftjTop� WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxFtpForcePasvIpComboLeftjTop� WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxFtpUseMlsdComboLeftjTop}WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  TEditFtpAccountEditLeft� TopWidthHeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrder TextFtpAccountEditOnChange
DataChange  	TComboBoxFtpHostComboLeftjTop� WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TCheckBoxVMSAllRevisionsCheckLeftTop� Width�HeightCaption(   Visa alla fil&revisioner på VMS-servrarTabOrder    	TTabSheetS3SheetTagHelpType	htKeywordHelpKeywordui_login_s3CaptionS3
ImageIndex
TabVisible
DesignSize��  	TGroupBoxS3GroupLeftTopWidth�HeighthAnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�h  TLabelLabel27Left	TopWidthNHeightCaption&Standardregion:FocusControlS3DefaultReqionCombo  TLabelS3UrlStyleLabelLeft	Top3Width3HeightCaption
&URL-stil:FocusControlS3UrlStyleCombo  	TComboBoxS3DefaultReqionComboLeft� TopWidthHeightAnchorsakLeftakTopakRight DropDownCount	MaxLength TabOrder TextS3DefaultRegionComboOnChange
DataChangeItems.Strings
af-south-1	ap-east-1	ap-east-2ap-northeast-1ap-northeast-2ap-northeast-3
ap-south-1
ap-south-2ap-southeast-1ap-southeast-2ap-southeast-3ap-southeast-4ap-southeast-5ap-southeast-7ca-central-1	ca-west-1
cn-north-1cn-northwest-1eu-central-1eu-central-2
eu-north-1
eu-south-1
eu-south-2	eu-west-1	eu-west-2	eu-west-3il-central-1me-central-1
me-south-1mx-central-1	sa-east-1	us-east-1	us-east-2us-gov-east-1us-gov-west-1	us-west-1	us-west-2   	TComboBoxS3UrlStyleComboLeft� Top0WidthHeightAutoCompleteStylecsDropDownListAnchorsakLeftakTopakRight 	MaxLength2TabOrderItems.Strings   Virtuell värd   Sökväg   	TCheckBoxS3RequesterPaysCheckLeftTopMWidth�HeightCaption   Begäranden &betalarTabOrder   	TGroupBoxS3AuthenticationGroupLeftToppWidth�Height� AnchorsakLeftakTopakRight CaptionAutentiseringTabOrder
DesignSize��   TLabelS3SessionTokenLabelLeft	TopWidthKHeightCaption&Sessionstoken:FocusControlS3SessionTokenMemo  TLabelS3RoleArnLabelLeft	Top� Width5HeightCaption
&Roll ARN:FocusControlS3RoleArnEdit  TMemoS3SessionTokenMemoLeft	Top$Width�Height]AnchorsakLeftakTopakRight 	MaxLength'TabOrder OnChange
DataChange	OnKeyDownNoteMemoKeyDown  TEditS3RoleArnEditLeft	Top� Width�HeightAnchorsakLeftakTopakRight TabOrderTextS3RoleArnEditOnChange
DataChange    	TTabSheetWebDavSheetTagHelpType	htKeywordHelpKeywordui_login_webdavCaptionWebDAV
ImageIndex
TabVisible
DesignSize��  	TGroupBoxWebdavGroupLeftTopWidth�Height1AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�1  	TCheckBoxWebDavLiberalEscapingCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption-&Tolerera icke-kodade specialtecken i filnamnTabOrder OnClick
DataChange    	TTabSheet	ConnSheetTagHelpType	htKeywordHelpKeywordui_login_connectionCaption
Anslutning
ImageIndex
TabVisible
DesignSize��  	TGroupBoxFtpPingGroupLeftTop� Width�Height|AnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSize�|  TLabelFtpPingIntervalLabelLeft	Top^Width� HeightCaptionSekunder &mellan keepalivesFocusControlFtpPingIntervalSecEdit  TUpDownEditFtpPingIntervalSecEditLeft Top[WidthPHeight	AlignmenttaRightJustifyMaxValue       �
@MinValue       ��?AnchorsakTopakRight 	MaxLengthTabOrderOnChange
DataChange  TRadioButtonFtpPingOffButtonLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption&AvTabOrder OnClick
DataChange  TRadioButtonFtpPingDummyCommandButtonLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption#   Kör kommandon för &dummy-protkollTabOrderOnClick
DataChange  TRadioButtonFtpPingDirectoryListingButtonLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption)   &Och läs dessutom den aktuella katalogenTabOrderOnClick
DataChange   	TGroupBoxTimeoutGroupLeftTopQWidth�Height4AnchorsakLeftakTopakRight Caption	TimeouterTabOrder
DesignSize�4  TLabelLabel11Left	TopWidth� HeightCaption   Timeout för se&rversvar:FocusControlTimeoutEdit  TLabelLabel12LeftvTopWidth+HeightAnchorsakTopakRight CaptionsekunderFocusControlTimeoutEdit  TUpDownEditTimeoutEditLeft TopWidthPHeight	AlignmenttaRightJustify	Increment       �@MaxValue      ��@MinValue       �@AnchorsakTopakRight 	MaxLengthTabOrder OnChange
DataChange   	TGroupBox	PingGroupLeftTop� Width�Height|AnchorsakLeftakTopakRight Caption
KeepalivesTabOrder
DesignSize�|  TLabelPingIntervalLabelLeft	Top^Width� HeightCaptionSekunder &mellan keepalivesFocusControlPingIntervalSecEdit  TUpDownEditPingIntervalSecEditLeft Top[WidthPHeight	AlignmenttaRightJustifyMaxValue       �
@MinValue       ��?AnchorsakTopakRight 	MaxLengthTabOrderOnChange
DataChange  TRadioButtonPingOffButtonLeftTopWidth�HeightAnchorsakLeftakTopakRight CaptionA&vTabOrder OnClick
DataChange  TRadioButtonPingNullPacketButtonLeftTop-Width�HeightAnchorsakLeftakTopakRight CaptionSkicka SSH-&null-paketTabOrderOnClick
DataChange  TRadioButtonPingDummyCommandButtonLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption%   Kör kommandon för &dummy-protokoll:TabOrderOnClick
DataChange   	TGroupBoxIPvGroupLeftTopWidth�Height1AnchorsakLeftakTopakRight Caption   Version för internetprotokollTabOrder TRadioButtonIPAutoButtonLeftTopWidtheHeightCaptionA&utomatiskTabOrder OnClick
DataChange  TRadioButton
IPv4ButtonLeft� TopWidtheHeightCaptionIPv&4TabOrderOnClick
DataChange  TRadioButton
IPv6ButtonLeft� TopWidtheHeightCaptionIPv&6TabOrderOnClick
DataChange   	TGroupBoxConnectionGroupLeftTopWidth�HeightIAnchorsakLeftakTopakRight Caption
AnslutningTabOrder 
DesignSize�I  	TCheckBoxFtpPasvModeCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   &Passivt lägeTabOrder OnClick
DataChange  	TCheckBoxBufferSizeCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption(   Optimera storlek på anslutnings&buffertTabOrderOnClick
DataChange    	TTabSheet
ProxySheetTagHelpType	htKeywordHelpKeywordui_login_proxyCaptionProxy
ImageIndex
TabVisible
DesignSize��  	TGroupBoxProxyTypeGroupLeftTopWidth�Height� AnchorsakLeftakTopakRight CaptionProxyTabOrder 
DesignSize��   TLabelProxyMethodLabelLeft	TopWidth:HeightCaption&Typ av proxy:FocusControlSshProxyMethodCombo  TLabelProxyHostLabelLeft	Top0Width[HeightCaption   Pro&xyns värdnamn:FocusControlProxyHostEdit  TLabelProxyPortLabelLeftGTop0WidthFHeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlProxyPortEdit  TLabelProxyUsernameLabelLeft	Top_Width;HeightCaption   &Användarnamn:FocusControlProxyUsernameEdit  TLabelProxyPasswordLabelLeft� Top_Width5HeightCaption   &Lösenord:FocusControlProxyPasswordEdit  	TComboBoxSshProxyMethodComboLeft� TopWidthyHeightStylecsDropDownListTabOrder OnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTPTelnetLokal   TUpDownEditProxyPortEditLeftGTopBWidthfHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrderOnChange
DataChange  TEditProxyHostEditLeft	TopBWidth8HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderTextProxyHostEditOnChange
DataChange  TEditProxyUsernameEditLeft	TopqWidth� Height	MaxLengthdTabOrderTextProxyUsernameEditOnChange
DataChange  TPasswordEditProxyPasswordEditLeft� TopqWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextProxyPasswordEditOnChange
DataChange  	TComboBoxFtpProxyMethodComboLeft� TopWidth!HeightStylecsDropDownListAnchorsakLeftakTopakRight DropDownCountTabOrderOnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTP
SITE %host!USER %proxyuser, USER %user@%host
OPEN %hostUSER %proxyuser, USER %userUSER %user@%hostUSER %proxyuser@%hostUSER %user@%host %proxyuserUSER %user@%proxyuser@%host   	TComboBoxNeonProxyMethodComboLeft� TopWidthyHeightStylecsDropDownListTabOrderOnChange
DataChangeItems.StringsIngenSOCKS4SOCKS5HTTP   TButtonProxyAutodetectButtonLeft	Top� WidthdHeightCaption&Automatisk identifieringTabOrderOnClickProxyAutodetectButtonClick   	TGroupBoxProxySettingsGroupLeftTop� Width�Height� AnchorsakLeftakTopakRight Caption   Inställningar proxyTabOrder
DesignSize��   TLabelProxyTelnetCommandLabelLeft	TopWidth]HeightCaptionTelnetko&mmando:FocusControlProxyTelnetCommandEdit  TLabelLabel17Left	TophWidth� HeightCaption-   Låt &DNS-namnuppslagningar göras av proxyn:FocusControlProxyDNSCombo  TLabelProxyLocalCommandLabelLeft	TopWidthyHeightCaptionLokalt proxyko&mmando:FocusControlProxyLocalCommandEdit  TEditProxyTelnetCommandEditLeft	Top(Width�HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextProxyTelnetCommandEditOnChange
DataChange  	TCheckBoxProxyLocalhostCheckLeftTopNWidth�HeightAnchorsakLeftakTopakRight Caption(   Låt lokala a&nslutningar gå via proxynTabOrder  	TComboBoxProxyDNSComboLeftjTopeWidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderItems.Strings
AutomatiskNejJa   TEditProxyLocalCommandEditLeft	Top(WidthLHeightAnchorsakLeftakTopakRight TabOrderTextProxyLocalCommandEditOnChange
DataChange  TButtonProxyLocalCommandBrowseButtonLeft[Top'WidthRHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClick"ProxyLocalCommandBrowseButtonClick  TStaticTextProxyTelnetCommandHintTextLeft^Top?WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption   mönsterTabOrderTabStop	  TStaticTextProxyLocalCommandHintTextLeftTop?WidthOHeight	AlignmenttaRightJustifyAnchorsakTopakRight AutoSizeCaption   mönsterTabOrderTabStop	    	TTabSheetTunnelSheetTagHelpType	htKeywordHelpKeywordui_login_tunnelCaptionTunnel
ImageIndex
TabVisible
DesignSize��  	TGroupBoxTunnelSessionGroupLeftTopWidth�HeightxAnchorsakLeftakTopakRight Caption    Värd för att sätta upp tunnelTabOrder
DesignSize�x  TLabelLabel6Left	TopWidth=HeightCaption   &Värdnamn:FocusControlTunnelHostNameEdit  TLabelLabel14LeftGTopWidthFHeightAnchorsakTopakRight CaptionPo&rtnummer:FocusControlTunnelPortNumberEdit  TLabelLabel15Left	TopEWidth;HeightCaption   &Användarnamn:FocusControlTunnelUserNameEdit  TLabelLabel16Left� TopEWidth5HeightCaption   &Lösenord:FocusControlTunnelPasswordEdit  TEditTunnelHostNameEditLeft	Top(Width8HeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder TextTunnelHostNameEditOnChange
DataChange  TEditTunnelUserNameEditLeft	TopWWidth� Height	MaxLengthdTabOrderTextTunnelUserNameEditOnChange
DataChange  TPasswordEditTunnelPasswordEditLeft� TopWWidth� HeightAnchorsakLeftakTopakRight 	MaxLengthdTabOrderTextTunnelPasswordEditOnChange
DataChange  TUpDownEditTunnelPortNumberEditLeftGTop(WidthfHeight	AlignmenttaRightJustifyMaxValue      ��@MinValue       ��?AnchorsakTopakRight TabOrderOnChange
DataChange   	TCheckBoxTunnelCheckLeft
TopWidth�HeightAnchorsakLeftakTopakRight CaptionAnslut med SSH-tunnelTabOrder OnClick
DataChange  	TGroupBoxTunnelOptionsGroupLeftTop� Width�Height4AnchorsakLeftakTopakRight Caption   Alternativ för tunnelTabOrder
DesignSize�4  TLabelLabel21Left	TopWidth]HeightCaption&Lokal tunnelport:FocusControlTunnelLocalPortNumberEdit  	TComboBoxTunnelLocalPortNumberEditLeftGTopWidthfHeightAutoCompleteAnchorsakTopakRight 	MaxLength2TabOrder TextTunnelLocalPortNumberEditOnChange
DataChangeItems.Strings   Välj automatiskt    	TGroupBoxTunnelAuthenticationParamsGroupLeftTop� Width�HeightGAnchorsakLeftakTopakRight CaptionTunnelautentiseringsparametrarTabOrder
DesignSize�G  TLabelLabel18Left	TopWidthOHeightCaptionPrivat nyc&kelfilFocusControlTunnelPrivateKeyEdit3  TFilenameEditTunnelPrivateKeyEdit3Left	Top(Width�HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEdit3AfterDialogFilter�PuTTY privata nyckelfiler (*.ppk)|*.ppk|Alla privata nyckelfiler (*.ppk;*.pem;*.key;id_*)|*.ppk;*.pem;*.key;id_*|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj privat nyckelfilClickKey@AnchorsakLeftakTopakRight TabOrder TextTunnelPrivateKeyEdit3OnChange
DataChange    	TTabSheetSslSheetTagHelpType	htKeywordHelpKeywordui_login_tlsCaptionTLS/SSL
ImageIndex
TabVisible
DesignSize��  	TGroupBoxTlsGroupLeftTopWidth�HeighthAnchorsakLeftakTopakRight CaptionTLS-alternativTabOrder 
DesignSize�h  TLabelMinTlsVersionLabelLeft	TopWidthwHeightCaptionMi&nimum TLS-version:FocusControlMinTlsVersionCombo  TLabelMaxTlsVersionLabelLeft	Top3WidthxHeightCaptionMa&ximal TLS-version:FocusControlMaxTlsVersionCombo  	TComboBoxMinTlsVersionComboLeftYTopWidthTHeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChangeMinTlsVersionComboChangeItems.StringsTLS 1.0TLS 1.1TLS 1.2TLS 1.3   	TComboBoxMaxTlsVersionComboLeftYTop0WidthTHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChangeMaxTlsVersionComboChangeItems.StringsTLS 1.0TLS 1.1TLS 1.2TLS 1.3   	TCheckBoxSslSessionReuseCheck2LeftTopMWidth�HeightAnchorsakLeftakTopakRight Caption3   Å&teranvänd TLS-sessions-ID för dataanslutningarTabOrderOnClick
DataChange   	TGroupBoxTlsAuthenticationGroupLeft	ToppWidth�HeightIAnchorsakLeftakTopakRight CaptionParametrar autentiseringTabOrder
DesignSize�I  TLabelLabel4Left	TopWidthlHeightCaptionKlientcertifikatfil:FocusControlTlsCertificateFileEdit  TFilenameEditTlsCertificateFileEditLeft	Top(Width�HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialog!TlsCertificateFileEditAfterDialogFilteriCertifikat och privata nyckelfiler (*.pfx;*.p12;*.key;*.pem)|*.pfx;*.p12;*.key;*.pem|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj klientcertifikatfilenClickKey@AnchorsakLeftakTopakRight TabOrder TextTlsCertificateFileEditOnChange
DataChange    	TTabSheetAdvancedSheetTagHelpType	htKeywordHelpKeywordui_login_sshCaptionSSH
ImageIndex
TabVisible
DesignSize��  	TGroupBoxProtocolGroupLeftTopWidth�Height1AnchorsakLeftakTopakRight Caption   Alternativ för protokollTabOrder 
DesignSize�1  	TCheckBoxCompressionCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Använd &komprimeringTabOrder OnClick
DataChange   	TGroupBoxEncryptionGroupLeftTop9Width�Height� AnchorsakLeftakTopakRight Caption   KrypteringsinställningarTabOrder
DesignSize��   TLabelLabel8Left	TopWidth� HeightCaption$   &Riktlinjer för krypteringschiffer:FocusControlCipherListBox  TListBoxCipherListBoxLeft	Top(WidthNHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  	TCheckBoxSsh2LegacyDESCheckLeftTop� Width�HeightAnchorsakLeftakRightakBottom Caption-   Tillåt arvsanvänding av single-&DES i SSH-2TabOrder  TButtonCipherUpButtonLeft]Top(WidthPHeightAnchorsakTopakRight Caption&UppTabOrderOnClickCipherButtonClick  TButtonCipherDownButtonLeft]TopGWidthPHeightAnchorsakTopakRight Caption&NerTabOrderOnClickCipherButtonClick    	TTabSheetKexSheetTagHelpType	htKeywordHelpKeywordui_login_kexCaption
Nyckelbyte
ImageIndex
TabVisible
DesignSize��  	TGroupBoxKexOptionsGroupLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption%   Alternativ för nyckelbytesalgoritmenTabOrder 
DesignSize�  TLabelLabel28Left	TopWidth� HeightCaption   Ri&ktlinjer för algoritmen:FocusControl
KexListBox  TListBox
KexListBoxLeft	Top(WidthNHeight� AnchorsakLeftakTopakRightakBottom DragModedmAutomatic
ItemHeightTabOrder OnClick
DataChange
OnDragDropAlgListBoxDragDrop
OnDragOverAlgListBoxDragOverOnStartDragAlgListBoxStartDrag  TButtonKexUpButtonLeft]Top(WidthPHeightAnchorsakTopakRight Caption&UppTabOrderOnClickKexButtonClick  TButtonKexDownButtonLeft]TopDWidthPHeightAnchorsakTopakRight Caption&NerTabOrderOnClickKexButtonClick  	TCheckBoxAuthGSSAPIKEXCheckLeftTop� WidthHeightAnchorsakLeftakBottom Caption!   Försök med &GSSAPI-nyckelutbyteTabOrderOnClick
DataChange   	TGroupBoxKexReexchangeGroupLeftTop Width�HeightQAnchorsakLeftakTopakRight Caption(   Alternativ för kontroll av nyckelutbyteTabOrder
DesignSize�Q  TLabelLabel31Left	TopWidth� HeightCaption?   Max antal minuter innan nyckeluppdatering (0 ger ingen gräns):Color	clBtnFaceFocusControlRekeyTimeEditParentColor  TLabelLabel32Left	Top3Width� HeightCaption<   Max antal data innan nyckeluppdatering (0 ger ingen gräns):Color	clBtnFaceFocusControlRekeyDataEditParentColor  TUpDownEditRekeyTimeEditLeft]TopWidthPHeight	AlignmenttaRightJustifyMaxValue       �	@AnchorsakTopakRight 	MaxLengthTabOrder OnChange
DataChange  TEditRekeyDataEditLeft]Top0WidthPHeightAnchorsakTopakRight 	MaxLength
TabOrderOnChange
DataChange    	TTabSheet	AuthSheetTagHelpType	htKeywordHelpKeywordui_login_authenticationCaptionAutentisering
ImageIndex

TabVisible
DesignSize��  	TCheckBoxSshNoUserAuthCheckLeft
TopWidth�HeightAnchorsakLeftakTopakRight Caption/   Kringgå autentisering helt och hållet (SSH-2)TabOrder OnClick
DataChange  	TGroupBoxAuthenticationGroupLeftTopWidth�Height_AnchorsakLeftakTopakRight Caption   Alternativ för autentiseringTabOrder
DesignSize�_  	TCheckBoxTryAgentCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption,   Försök använda autentisering med &PageantTabOrder OnClick
DataChange  	TCheckBoxAuthKICheckLeftTop-Width�HeightAnchorsakLeftakTopakRight CaptionA   Försök använda 'tangentbords&interaktiv' autentisering (SSH-2)TabOrderOnClick
DataChange  	TCheckBoxAuthKIPasswordCheckLeftTopDWidth�HeightAnchorsakLeftakTopakRight Caption)   Svara med lösenord vid första &promptenTabOrderOnClick
DataChange   	TGroupBoxAuthenticationParamsGroupLeftTop~Width�Height� AnchorsakLeftakTopakRight CaptionParametrar autentiseringTabOrder
DesignSize��   TLabelPrivateKeyLabelLeft	Top-WidthOHeightCaptionPrivat nyc&kelfilFocusControlPrivateKeyEdit3  TLabelDetachedCertificateLabelLeft	TopyWidth� HeightCaption1   Certifikat att &använda med den privata nyckeln:FocusControlDetachedCertificateEdit  	TCheckBoxAgentFwdCheckLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Tillåt agent-vidarebe&fordranTabOrder OnClick
DataChange  TFilenameEditPrivateKeyEdit3Left	Top?Width�HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEdit3AfterDialogFilter�PuTTY privata nyckelfiler (*.ppk)|*.ppk|Alla privata nyckelfiler (*.ppk;*.pem;*.key;id_*)|*.ppk;*.pem;*.key;id_*|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj privat nyckelfilClickKey@AnchorsakLeftakTopakRight TabOrderTextPrivateKeyEdit3OnChange
DataChange  TButtonPrivateKeyToolsButtonLeft� TopZWidth^HeightCaption&VerktygTabOrderOnClickPrivateKeyToolsButtonClick  TButtonPrivateKeyViewButtonLeft	TopZWidth� HeightCaption&Visa publik nyckelTabOrderOnClickPrivateKeyViewButtonClick  TFilenameEditDetachedCertificateEditLeft	Top� Width�HeightAcceptFiles	OnBeforeDialogPathEditBeforeDialogOnAfterDialogPrivateKeyEdit3AfterDialogFilter5Public nyckelfiler (*.pub)|*.pub|Alla filer (*.*)|*.*DialogOptions
ofReadOnlyofPathMustExistofFileMustExist DialogTitle   Välj certifikatfilClickKey@AnchorsakLeftakTopakRight TabOrderTextDetachedCertificateEditOnChange
DataChange   	TGroupBoxGSSAPIGroupLeftTop0Width�HeightHAnchorsakLeftakTopakRight CaptionGSSAPITabOrder
DesignSize�H  	TCheckBoxAuthGSSAPICheck3LeftTopWidth�HeightAnchorsakLeftakTopakRight Caption3   Försök använda GSSAPI/SSPI autentisering (SSH-2)TabOrder OnClickAuthGSSAPICheck3Click  	TCheckBoxGSSAPIFwdTGTCheckLeftTop-Width�HeightAnchorsakLeftakTopakRight Caption4   Tillåt GSSAPI &vidarbefodra autentiseringsuppgifterTabOrderOnClickAuthGSSAPICheck3Click    	TTabSheet	BugsSheetTagHelpType	htKeywordHelpKeywordui_login_bugsCaptionBuggar
ImageIndex	
TabVisible
DesignSize��  	TGroupBoxBugsGroupBoxLeftTopWidth�HeightAnchorsakLeftakTopakRight Caption   Upptäcka buggar i SSH-servrarTabOrder 
DesignSize�  TLabelBugHMAC2LabelLeft	TopPWidth� HeightCaption(   Beräkningsfel av H&MAC-nycklar i SSH-2:FocusControlBugHMAC2Combo  TLabelBugDeriveKey2LabelLeft	TopmWidth� HeightCaption.   Beräkningsf&el av krypteringsnycklar i SSH-2:FocusControlBugDeriveKey2Combo  TLabelBugRSAPad2LabelLeft	Top� Width� HeightCaption-   Kräver &utfyllnad av RSA-signaturer i SSH-2:FocusControlBugRSAPad2Combo  TLabelBugPKSessID2LabelLeft	Top� Width� HeightCaption1Sessio&ns-id i SSH-2 PK autentisering missbrukas:FocusControlBugPKSessID2Combo  TLabelBugRekey2LabelLeft	Top� Width� HeightCaption%   Hanterar SSH-2 nyc&kelutbyte dåligt:FocusControlBugRekey2Combo  TLabelBugMaxPkt2LabelLeft	Top� Width� HeightCaption+   Ignorerar SSH-2 ma&ximum för paketstorlek:FocusControlBugMaxPkt2Combo  TLabelBugIgnore2LabelLeft	TopWidth� HeightCaption(Stannar vid ignore-meddelanden i SSH-&2:FocusControlBugIgnore2Combo  TLabelBugWinAdjLabelLeft	Top3Width� HeightCaption,   Stannar på WinSCP:s SSH-2 'winadj' begäranFocusControlBugWinAdjCombo  	TComboBoxBugHMAC2ComboLeftjTopMWidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugDeriveKey2ComboLeftjTopjWidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugRSAPad2ComboLeftjTop� WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugPKSessID2ComboLeftjTop� WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugRekey2ComboLeftjTop� WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugMaxPkt2ComboLeftjTop� WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange  	TComboBoxBugIgnore2ComboLeftjTopWidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrder OnChange
DataChange  	TComboBoxBugWinAdjComboLeftjTop0WidthCHeightStylecsDropDownListAnchorsakTopakRight TabOrderOnChange
DataChange    	TTabSheet	NoteSheetHelpType	htKeywordHelpKeywordui_login_noteCaption
Anteckning
ImageIndex
TabVisible
DesignSize��  	TGroupBox	NoteGroupLeftTopWidth�Height~AnchorsakLeftakTopakRightakBottom Caption
AnteckningTabOrder 
DesignSize�~  TMemoNoteMemoLeft	TopWidth�Height^AnchorsakLeftakTopakRightakBottom 	MaxLength�TabOrder OnChange
DataChange	OnKeyDownNoteMemoKeyDown     TPanel	LeftPanelLeft Top Width� Height�AlignalLeft
BevelOuterbvNoneTabOrder 
DesignSize� �  TPanelNavigationPanelLeftTopWidth� Height~AnchorsakLeftakTopakRightakBottom 
BevelOuterbvNoneTabOrder  	TTreeViewNavigationTreeLeft Top Width� Height~AlignalClientDoubleBuffered	HideSelectionHotTrack	IndentParentDoubleBufferedReadOnly	ShowButtonsShowRootTabOrder OnChangeNavigationTreeChangeOnCollapsingNavigationTreeCollapsingItems.NodeData
W     6               ����           E n v i r o n m e n t X 6               ����            D i r e c t o r i e s X 6               ����            R e c y c l e   b i n X 4           ��������            E n c r y p t i o n X (               ����            S F T P X &               ����            S C P X &           ��������            F T P X $               ����            S 3 X ,           ��������            W e b D A V X 4               ����           C o n n e c t i o n X *               ����            P r o x y X ,               ����            T u n n e l X &               ����           S S H X 8               ����            K e x   e x c h a n g e X <               ����            A u t h e n t i c a t i o n X (               ����            B u g s X (               ����            N o t e X      TButtonOKBtnLeftgTop�WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButton	CancelBtnLeft�Top�WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftTop�WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonColorButtonLeftTop�WidthPHeightAnchorsakLeftakBottom Caption   &FärgTabOrderOnClickColorButtonClick  
TImageListColorImageListAllocByLeft$Top!Bitmap
&  IL  P   �������������BM6       6   (   @                                                                                                                                                                                                                                                                                                                K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5                                                                                                                                                                                                                                         K?5 K?5 K?5 K?5                                                                                                                                                                                                                             dYQ K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                         K?5 s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R s`R K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         K?5 � � � � � � � � � � � � K?5                                                                                                                                                                                                         bXO K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   @            �                       ��� ��      �      �?      �      �      �      �      �      �      �      �      �      �      �      ��      ��                              
TImageListColorImageList120AllocByHeightWidthLeft� Top!Bitmap
�  IL     �������������BM6       6   (   P                                                                                                                                                                                                                                                                                                                                                                                    bXO K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                         K?5 ��o ��o ��o ��o ��o ��o ��o ��o K?5                                                                                                                                                                                                                                                                                         bXO K?5 K?5 0(" 0(" 0(" 0(" K?5 K?5 bXO                                                                                                                                                                                                                                                                                                     '! '! '! '!                                                                                                                                                                                                                                                                                     qg_ K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 qg_                                                                                                                                                                                                                                                         K?5 ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x )�> )�> ��x K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         K?5 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � K?5                                                                                                                                                                                                                                                         oe] K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 oe]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   P            �                       ��� ���         ��         ��         ��         ��         �          �          �          �          �          �          �          �          �          �          �          �          �          ���         ���                                 
TImageListColorImageList144AllocByHeightWidthLeft$TopQBitmap
�%  IL h t   �������������BM6       6   (   `              $                                                                                                                                                                                                                                                                                                                                                                                                                                          bXO K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                                                                                 K?5 ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o K?5                                                                                                                                                                                                                                                                                                                                                 K?5 s`R s`R s`R K?5 K?5 K?5 K?5 s`R s`R s`R K?5                                                                                                                                                                                                                                                                                                                                                 bXO K?5 K?5 K?5 B7/ B7/ B7/ B7/ K?5 K?5 K?5 bXO                                                                                                                                                                                                                                                                                                                                                                 0(" 0(" 0(" 0("                                                                                                                                                                                                                                                                                                                                             tjc K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 tjc                                                                                                                                                                                                                                                                                                         K?5 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 NB8 )�> )�> NB8 K?5                                                                                                                                                                                                                                                                                                         K?5 QD; ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x QD; K?5                                                                                                                                                                                                                                                                                                         K?5 UG= � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � UG= K?5                                                                                                                                                                                                                                                                                                         K?5 XJ? � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � XJ? K?5                                                                                                                                                                                                                                                                                                         K?5 [MB � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � [MB K?5                                                                                                                                                                                                                                                                                                         K?5 ^PD � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ^PD K?5                                                                                                                                                                                                                                                                                                         K?5 bSG � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � bSG K?5                                                                                                                                                                                                                                                                                                         K?5 eUI � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � eUI K?5                                                                                                                                                                                                                                                                                                         K?5 iXL � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � iXL K?5                                                                                                                                                                                                                                                                                                         K?5 l[N � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � l[N K?5                                                                                                                                                                                                                                                                                                         K?5 o^Q � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � o^Q K?5                                                                                                                                                                                                                                                                                                         K?5 saS � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � saS K?5                                                                                                                                                                                                                                                                                                         K?5 vdV � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � vdV K?5                                                                                                                                                                                                                                                                                                         K?5 yfX �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g �]g yfX K?5                                                                                                                                                                                                                                                                                                         ria OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 OC8 ria                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BM>       >   (   `                                   ��� ���         � ?         � ?         � ?         � ?         ���         �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          ���         ���                                 
TImageListColorImageList192AllocByHeight Width Left� TopQBitmap
�B  IL ` l     �������������BM6       6   (   �               @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  i_W K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 i_W                                                                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o ��o K?5                                                                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 s`R s`R s`R s`R K?5 K?5 K?5 K?5 K?5 K?5 s`R s`R s`R s`R K?5                                                                                                                                                                                                                                                                                                                                                                                                                                                                 i_W K?5 K?5 K?5 K?5 E:1 E:1 E:1 E:1 E:1 E:1 K?5 K?5 K?5 K?5 i_W                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     90( 90( 90( 90( 90( 90(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         -&  -&  -&  -&  -&  -&                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��~ L@6 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 L@6 ���                                                                                                                                                                                                                                                                                                                                                                                                                 L@6 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 MA8 L@6                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: PC: )�> )�> )�> PC: K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 RE; ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x ��x RE; K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 TG= � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � TG= K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 WI? � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � WI? K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 YK@ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � YK@ K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 [MB � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � [MB K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 ^OD � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ^OD K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 `QF � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � `QF K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 bSG � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � bSG K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 eUI � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � eUI K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 gWK � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � gWK K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 jYL � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � jYL K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 l[N � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � l[N K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 o]P � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � o]P K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 q_R � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � q_R K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 saS � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � saS K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 ucU � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ucU K?5                                                                                                                                                                                                                                                                                                                                                                                                                 K?5 xeW � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � xeW K?5                                                                                                                                                                                                                                                                                                                                                                                                                 L@6 zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY zgY L@6                                                                                                                                                                                                                                                                                                                                                                                                                 ��} K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 K?5 L@6 ��~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         BM>       >   (   �                                    ��� ����            ����            �  �            �  �            �  �            �  �            ���            ���            �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              �              ����            ����                                    
TPopupMenuPrivateKeyMenuLeft� Top� 	TMenuItemPrivateKeyGenerateItemCaption(&Generera nytt nyckelpar med PuTTYgen...OnClickPrivateKeyGenerateItemClick  	TMenuItemPrivateKeyUploadItemCaption%&Installera publik nyckel i server...OnClickPrivateKeyUploadItemClick       TPF0TSymlinkDialogSymlinkDialogLeft�Top� HelpType	htKeywordHelpKeyword
ui_symlinkBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSymlinkDialogClientHeight� ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenterOnShowFormShow
DesignSize��  
TextHeight 	TGroupBoxSymlinkGroupLeftTopWidth�Height� AnchorsakLeftakTopakRightakBottom TabOrder 
DesignSize��   TLabelFileNameLabelLeft	Top	Width]HeightCaption   &Länk/genväg fil:FocusControlFileNameEdit  TLabelLabel1Left	Top8WidthtHeightCaption   &Pekar länk/genväg till:FocusControlPointToEdit  TEditFileNameEditLeft	TopWidthHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrder OnChangeControlChange  TEditPointToEditLeft	TopJWidthHeightAnchorsakLeftakTopakRight 	MaxLength� TabOrderOnChangeControlChange  	TCheckBoxHardLinkCheckLeftTopgWidth�HeightCaption   &Hård länkTabOrderOnClickControlChange   TButtonOkButtonLeft� Top� WidthPHeightAnchorsakRightakBottom CaptionOKDefault	ModalResultTabOrder  TButtonCancelButtonLeft� Top� WidthPHeightAnchorsakRightakBottom Cancel	CaptionAvbrytModalResultTabOrder  TButton
HelpButtonLeftITop� WidthPHeightAnchorsakRightakBottom Caption   &HjälpTabOrderOnClickHelpButtonClick   TPF0TSynchronizeChecklistDialogSynchronizeChecklistDialogLeft4Top� HelpType	htKeywordHelpKeywordui_synchronize_checklistBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp CaptionSynchronization checklist XClientHeight	ClientWidth�Color	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 	Icon.Data
��      @@     (B  v   00     �%  �B  ((     h  Fh         �  ��       �	  V�       �  ޜ       h  ��  (   @   �           B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           p�K p�� p�� o�� o�� o�� n�� n�� m�� m�� m�� l�� l�� l�� k�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� i�K                                                                                 p�� p�� p�� p�� o�� o�� o�� n�� n�� n�� m�� m�� m�� l�� l�� l�� k�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                                                 q�� q�� q�� p�� p�� p�� o�� o�� o�� n�� n�� m�� m�� m�� l�� l�� l�� k�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                                                 r�� r�� q�� q�� p�� p�� p�� o�� o�� o�� n�� n�� n�� m�� m�� m�� l�� l�� l�� k�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                                                 r�� r�� r�� q�� q�� q�� p�� p�� p�� o�� o�� o�� n�� n�� m�� m�� m�� l�� l�� l�� k�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                                                 s�� s�� r�� r�� r�� q�� q�� p�� p�� p�� o�� o�� o�� n�� n�� n�� m�� m�� m�� l�� l�� l�� k�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                                                 s�� s�� s�� r�� r�� r���������������������������������������������������������������������������������������������������������������������������������� j�� j�� j�� j�� j�� j��                                                                                 t�� t�� s�� s�� s�� r���������������������������������������������������������������������������������������������������������������������������������� j�� j�� j�� j�� j�� j��                                                                                 t�� t�� t�� s�� s�� s���������������������������������������������������������������������������������������������������������������������������������� j�� j�� j�� j�� j�� j��                                                                                 u�� u�� t�� t�� t�� s���������������������������������������������������������������������������������������������������������������������������������� j�� j�� j�� j�� j�� j��                                                                                 v�� u�� u�� t�� t�� t��������������������������������������������������Ku��1`�������������������������������������������������������������������������� j�� j�� j�� j�� j�� j��                                                                                 v�� v�� u�� u�� u�� t����������������������������������������������4c��=��=��@l���������������������������������������������������������������������� j�� j�� j�� j�� j�� j��                                                                                 v�� v�� v�� v�� u�� u������������������������������������������Al��=��=��=��=���������������������������������������������������������������������� j�� j�� j�� j�� j�� j��                                                                                 w�� w�� v�� v�� v�� u��������������������������������������Ox��=��=��=��=��=�� S������������������������������������������������������������������ j�� j�� j�� j�� j�� j��                                                                                 x�� w�� w�� v�� v�� v����������������������������������]���=��=��>������)Z��=��=������������������������������������������������������������������ j�� j�� j�� j�� j�� j��                                                                                 x�� x�� w�� w�� w�� v������������������������������o���=��=��=��������������=��=��F�������������������������������������������������������������� k�� k�� j�� j�� j�� j��                                                                                 y�� x�� x�� x�� w�� w������������������������������=��=��=������������������Lu��=��=��]����������������������������������������������������������� k�� k�� k�� j�� j�� j��                                                                                 y�� y�� y�� x�� x�� w��������������������������=��=��=��y�����������������������A��=��=���������������������������������������������������������� l�� l�� k�� k�� k�� j��                                                                                 z�� y�� y�� y�� x�� x����������������������>��=��=��e���������������������������u���=��=��3b������������������������������������������������������ l�� l�� l�� k�� k�� k��                                                                                 z�� z�� y�� y�� y�� y������������������A��=��=��W}����������������������������������M��=��=������������������������������������������������������ m�� m�� l�� l�� l�� k��                                                                                 {�� z�� z�� z�� y�� y��������������L��=��=��Is������������������������������������������=��=��M�������������������������������������������������� m�� m�� m�� l�� l�� l��                                                                                 {�� {�� {�� z�� z�� y��������������-]��=��;h����������������������������������������������5c��=��=��s����������������������������������������������� n�� n�� m�� m�� m�� l��                                                                                 |�� {�� {�� {�� z�� z��������������������������������������������������������������������������>��=��A���������������������������������������������� o�� n�� n�� m�� m�� m��                                                                                 |�� |�� |�� {�� {�� {��������������������������������������������������������������������������]���=��=��Lu������������������������������������������ o�� o�� n�� n�� n�� m��                                                                                 }�� |�� |�� |�� {�� {������������������������������������������������������������������������������F��=��=������������������������������������������ p�� o�� o�� o�� n�� n��                                                                                 }�� }�� }�� |�� |�� |����������������������������������������������������������������������������������=��=��'Y�������������������������������������� p�� p�� o�� o�� o�� n��                                                                                 ~�� }�� }�� }�� |�� |����������������������������������������������������������������������������������"U��=��=�������������������������������������� q�� p�� p�� p�� o�� o��                                                                                 ~�� ~�� ~�� }�� }�� }��������������������������������������������������������������������������������������=��=��I���������������������������������� q�� q�� p�� p�� p�� o��                                                                                 �� �� ~�� ~�� }�� }��������������������������������������������������������������������������������������Bm��=��=��g������������������������������� r�� q�� q�� q�� p�� p��                                                                                 �� �� �� ~�� ~�� ~������������������������������������������������������������������������������������������@��=��>������������������������������ r�� r�� r�� q�� q�� p��                                                                                 ��� ��� �� �� �� ~������������������������������������������������������������������������������������������i���=��=��>j�������������������������� s�� r�� r�� r�� q�� q��                                                                                 ��� ��� ��� �� �� ����������������������������������������������������������������������������������������������J��=��=�������������������������� s�� s�� s�� r�� r�� r��                                                                                 ��� ��� ��� ��� ��� ��������������������������������������������������������������������������������������������������=��=�� S���������������������� t�� s�� s�� s�� r�� r��                                                                                 ��� ��� ��� ��� ��� ���������������������������������������������������������������������������������������������������+\��=��=���������������������� t�� t�� t�� s�� s�� s��                                                                                 ��� ��� ��� ��� ��� �������������������������������������������������������������������������������������������������������=��=��D������������������ u�� t�� t�� t�� s�� s��                                                                                 ��� ��� ��� ��� ��� �������������������������������������������������������������������������������������������������������Px��=��=��Y�������������� u�� u�� u�� t�� t�� t��                                                                                 ��� ��� ��� ��� ��� �����������������������������������������������������������������������������������������������������������
C��=��I�������������� v�� v�� u�� u�� t�� t��                                                                                 ��� ��� ��� ��� ��� ���������������������������������������������������������������������������������������������������������������+\������������������ v�� v�� v�� u�� u�� u��                                                                                 ��� ��� ��� ��� ��� ����������������������������������������������������������������������������������������������������������������������������������� w�� v�� v�� v�� v�� u��                                                                                 ��� ��� ��� ��� ��� ����������������������������������������������������������������������������������������������������������������������������������� w�� w�� w�� v�� v�� v��                                                                                 ��� ��� ��� ��� ��� ����������������������������������������������������������������������������������������������������������������������������������� x�� x�� w�� w�� v�� v��                                                                                 ��� ��� ��� ��� ��� ����������������������������������������������������������������������������������������������������������������������������������� y�� x�� x�� w�� w�� w��                                                                                 ��� ��� ��� ��� ��� ����������������������������������������������������������������������������������������������������������������������������������� y�� y�� x�� x�� x�� w��                                                                                 ��� ��� ��� ��� ��� ����������������������������������������������������������������������������������������������������������������������������������� y�� y�� y�� y�� x�� x��                                                                                 ��� ��� ��� ��� ��� ��������������������������������������������������������������������������������������������������������������� z�� z�� y�� y�� y�� x��                                                                                 ��� ��� ��� ��� ��� ��������������������������������������������������������������������������������������������������������������� {�� z�� z�� y�� y�� y��                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���������j���i���h���g���f���e���d���c���b���b���a���`���_���^���]���\��������� j�� j�� |�� |�� |�� {�� {�� {�� z�� z�� z�� y��                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���������m���m���l���k���j���i���h���g���f���e���d���c���b���a���`���_��������� j�� j�� }�� }�� |�� |�� |�� {�� {�� {�� z�� z��                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���������q���p���o���n���m���l���k���j���i���h���g���g���f���e���d���c��������� j�� j�� }�� }�� }�� |�� |�� |�� {�� {�� {�� {��                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���������t���s���r���r���q���p���o���n���m���l���k���j���i���h���g���f��������� j�� j�� ~�� ~�� }�� }�� }�� |�� |�� |�� |�� ���                                                                                 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��������������������������������������������������������������� j�� v�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                 �ŀ ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��������������������������������������������������������������� v�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �À                                                                                                                                ��(��|������������������������������������������������|��&                                                                                                                                                                                            ��(��������������        ����������������&                                                                                                                                                                                                            ��������������        ��������������                                                                                                                                                                                                                ����������������������������������                                                                                                                                                                                                                ��k��������������������������������i                                                                                                                                                                                                                 �������������������������������� ��                                                                                                                                                                                                                    ����������������������������                                                                                                                                                                                                                             ����l��������������l ��                                                                                                                                                                                                                                                                                                                                                                                ��������������������������    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ���    ����  ?�������������������������������������������������������������(   0   `          �%                                                                                                                                                                                                                                                                                                                                                                                                                                               p�} p�� o�� o�� o�� n�� n�� m�� m�� l�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�}                                                         q�� q�� p�� p�� o�� o�� n�� n�� m�� m�� m�� l�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                         r�� q�� q�� p�� p�� o�� o�� o�� n�� n�� m�� m�� l�� l�� k�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                         r�� r�� q�� q�� q�� p�� p�� o�� o�� n�� n�� m�� m�� m�� l�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                         s�� s�� r�� r���������������������������������������������������������������������������������������������������������� j�� j�� j�� j��                                                         t�� s�� s�� r���������������������������������������������������������������������������������������������������������� j�� j�� j�� j��                                                         t�� t�� t�� s���������������������������������������������������������������������������������������������������������� j�� j�� j�� j��                                                         u�� u�� t�� t���������������������������������������������������������������������������������������������������������� j�� j�� j�� j��                                                         v�� u�� u�� t������������������������������������������
C��Al���������������������������������������������������������� j�� j�� j�� j��                                                         v�� v�� v�� u��������������������������������������
C��=��=���������������������������������������������������������� j�� j�� j�� j��                                                         w�� w�� v�� v����������������������������������F��=��	B��=��P������������������������������������������������������ j�� j�� j�� j��                                                         x�� w�� w�� v������������������������������L��=��$V������G��=��y��������������������������������������������������� j�� j�� j�� j��                                                         x�� x�� x�� w�������������������������� S��=��P��������������=��
C�������������������������������������������������� k�� k�� j�� j��                                                         y�� y�� x�� x����������������������,]��=��L������������������&X��=��Rz���������������������������������������������� l�� k�� k�� j��                                                         z�� y�� y�� y������������������6d��=��F��������������������������=��=���������������������������������������������� l�� l�� k�� k��                                                         {�� z�� z�� y��������������Lu��=��A������������������������������Jt��=��-]������������������������������������������ m�� m�� l�� l��                                                         {�� {�� z�� z��������������1`��@��������������������������������������@��=������������������������������������������ n�� m�� m�� l��                                                         |�� {�� {�� {����������������������������������������������������������s���=��J�������������������������������������� n�� n�� m�� m��                                                         }�� |�� |�� {��������������������������������������������������������������M��=��k����������������������������������� o�� o�� n�� n��                                                         }�� }�� |�� |������������������������������������������������������������������=��@���������������������������������� p�� o�� o�� n��                                                         ~�� }�� }�� }������������������������������������������������������������������1`��=��Bm������������������������������ p�� p�� p�� o��                                                         �� ~�� ~�� }����������������������������������������������������������������������=��=������������������������������ q�� q�� p�� p��                                                         �� �� ~�� ~����������������������������������������������������������������������W}��=��$V�������������������������� r�� q�� q�� p��                                                         ��� �� �� ��������������������������������������������������������������������������D��=�������������������������� r�� r�� r�� q��                                                         ��� ��� ��� ������������������������������������������������������������������������������=��F���������������������� s�� s�� r�� r��                                                         ��� ��� ��� ������������������������������������������������������������������������������� S��=��]������������������� t�� s�� s�� r��                                                         ��� ��� ��� �����������������������������������������������������������������������������������=��>������������������ t�� t�� t�� s��                                                         ��� ��� ��� �����������������������������������������������������������������������������������>j��=��=i�������������� u�� u�� t�� t��                                                         ��� ��� ��� ���������������������������������������������������������������������������������������D��Gq�������������� v�� u�� u�� t��                                                         ��� ��� ��� ����������������������������������������������������������������������������������������������������������� v�� v�� v�� u��                                                         ��� ��� ��� ����������������������������������������������������������������������������������������������������������� w�� w�� v�� v��                                                         ��� ��� ��� ����������������������������������������������������������������������������������������������������������� x�� w�� w�� v��                                                         ��� ��� ��� ����������������������������������������������������������������������������������������������������������� y�� x�� x�� w��                                                         ��� ��� ��� ����������������������������������������������������������������������������������������������������������� y�� y�� x�� x��                                                         ��� ��� ��� ��������������������������������������������������������������������������������������������� z�� y�� y�� y��                                                         ��� ��� ��� ������������������������������j���i���g���f���e���d���c���b���`���_���^���]������������������������������ {�� z�� z�� y��                                                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ������n���m���k���j���i���g���g���e���d���c���b���`������ j�� }�� }�� }�� |�� |�� {�� {�� z�� z��                                                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ������r���p���o���n���m���l���j���i���h���g���e���d������ j�� ~�� ~�� }�� }�� |�� |�� {�� {�� }��                                                         ��� ��� ��� ��� ��� ��� ��� ��� ��� ������K���K���J���J���I���H���H���G���F���E���E���D������ j�� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                         �Ŗ ��� ��� ��� ��� ��� ��� ��� ��� ��������������������������������������������� v�� ��� ��� ��� ��� ��� ��� ��� ��� �Ľ                                                                                                ��M������������������������������������E                                                                                                                                                ��_���������        ������������                                                                                                                                                        ��F�����������4��4�����������q                                                                                                                                                        ��
��������������������������                                                                                                                                                            ��W��������������������[                                                                                                                                                                    ��A��������������9                                                                                    ������  ������  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �����  �����  �����  �����  �����  �����  (   (   P          @                                                                                                                                                                                                                                                                                                                                                                           p�� p�� o�� o�� n�� n�� m�� m�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                 q�� q�� p�� p�� o�� n�� n�� m�� m�� l�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                 r�� r�� q�� p�� p�� o�� o�� n�� n�� m�� m�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                                 s�� r�� r������������������������������������������������������������������������������������������ j�� j�� j��                                                 t�� s�� s������������������������������������������������������������������������������������������ j�� j�� j��                                                 u�� t�� t������������������������������������������������������������������������������������������ j�� j�� j��                                                 u�� u�� t������������������������������������������������������������������������������������������ j�� j�� j��                                                 v�� v�� u����������������������������������A��=�������������������������������������������������� j�� j�� j��                                                 w�� w�� v������������������������������F��>��=��&X���������������������������������������������� j�� j�� j��                                                 x�� w�� w��������������������������J��=������Y��=���������������������������������������������� j�� j�� j��                                                 y�� x�� x����������������������O��=��������������D��F������������������������������������������ k�� k�� j��                                                 z�� y�� y������������������ S��=��q�������������������=��]��������������������������������������� l�� k�� k��                                                 {�� z�� y��������������,]��=��a����������������������� S��>�������������������������������������� m�� l�� l��                                                 {�� {�� z��������������=��Qy������������������������������=��7e���������������������������������� n�� m�� m��                                                 |�� |�� {��������������������������������������������������>j��=���������������������������������� o�� n�� m��                                                 }�� }�� |������������������������������������������������������>��O������������������������������ o�� o�� n��                                                 ~�� }�� }������������������������������������������������������g���=��w��������������������������� p�� p�� o��                                                 �� ~�� ~����������������������������������������������������������I��
C�������������������������� q�� q�� p��                                                 ��� �� ��������������������������������������������������������������=��Nw���������������������� r�� q�� q��                                                 ��� ��� ��������������������������������������������������������������'Y��=���������������������� s�� r�� r��                                                 ��� ��� �������������������������������������������������������������������=��+\������������������ t�� s�� s��                                                 ��� ��� �������������������������������������������������������������������Lu��=������������������ t�� t�� s��                                                 ��� ��� �����������������������������������������������������������������������A��J�������������� u�� u�� t��                                                 ��� ��� �����������������������������������������������������������������������w���A�������������� v�� v�� u��                                                 ��� ��� ������������������������������������������������������������������������������������������� w�� v�� v��                                                 ��� ��� ������������������������������������������������������������������������������������������� x�� w�� w��                                                 ��� ��� ������������������������������������������������������������������������������������������� y�� x�� x��                                                 ��� ��� ������������������������������������������������������������������������������������������� z�� y�� y��                                                 ��� ��� ������������������������������������������������������������������������������� z�� z�� y��                                                 ��� ��� ��� ��� ��� ��� ��� ������j���i���g���f���d���c���a���`���^���]������ j�� }�� }�� |�� |�� {�� {�� z��                                                 ��� ��� ��� ��� ��� ��� ��� ������o���m���l���j���i���g���f���d���c���b������ j�� ~�� ~�� }�� }�� |�� |�� {��                                                 ��� ��� ��� ��� ��� ��� ��� ������s���r���p���o���m���l���j���i���g���f������ j�� ��� ��� �� ~�� ~�� ~�� ���                                                 �ǵ ��� ��� ��� ��� ��� ��� ��������������������������������������� {�� ��� ��� ��� ��� ��� ��� �ǵ                                                     y� �� �� �� �� �� ����Y��������������Q��Q��������������Z �� �� �� �� �� �� y�                                                                                            ���������        ���������                                                                                                                                ������������������������                                                                                                                                ��&��������������������&                                                                                                                                    ��>��������������>                                                                    �����   �����   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �   ?   �      ����   �� ��   �� ��   �����   (       @          �                                                                                                                                                                                                                                                                                                       o�� p�� o�� n�� m�� m�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                         q�� q�� p�� o�� o�� n�� m�� l�� l�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                         r�� r�� q�� p�� p�� o�� n�� m�� m�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� j��                                         s�� s�� r������������������������������������������������������������������ j�� j�� j��                                         t�� t�� s������������������������������������������������������������������ j�� j�� j��                                         v�� u�� t��������������������������0`�������������������������������������� j�� j�� j��                                         w�� v�� u����������������������L��=��7e���������������������������������� j�� j�� j��                                         x�� w�� v������������������ S�� S������=���������������������������������� j�� j�� j��                                         y�� x�� w��������������,]��L����������Bm��P������������������������������ k�� k�� j��                                         z�� y�� x����������;h��F������������������@��{��������������������������� l�� l�� k��                                         {�� z�� y����������A����������������������k���
C�������������������������� m�� m�� l��                                         |�� {�� z��������������������������������������J��T{���������������������� o�� n�� m��                                         }�� |�� {������������������������������������������=���������������������� p�� o�� n��                                         ~�� }�� |������������������������������������������-]��-]������������������ q�� p�� o��                                         �� ~�� }����������������������������������������������=������������������ r�� q�� p��                                         ��� �� ����������������������������������������������Rz��J�������������� s�� r�� q��                                         ��� ��� ���������������������������������������������������
C��k����������� t�� s�� r��                                         ��� ��� ���������������������������������������������������y���@���������� u�� t�� s��                                         ��� ��� �������������������������������������������������������(Z���������� v�� u�� t��                                         ��� ��� ������������������������������������������������������������������� w�� v�� v��                                         ��� ��� ������������������������������������������������������������������� x�� w�� w��                                         ��� ��� ������������������������������������������������������������������� y�� x�� x��                                         ��� ��� ���������������)���(���,���,���,���,���,���,���,���,��������������� z�� y�� y��                                         ��� ��� ���������������d���b���`���^���\���[���Z���X������u�������� {�� z�� z��                                         ��� ��� ��� ��� ��� ������r���p���n���l���j���h���g���e������ j�� }�� }�� |�� {�� }��                                         ��� ��� ��� ��� ��� ������"���"���"���"���!���!���!���!������ v�� ��� ��� ��� ��� ���                                         �� ��, ��, ��, ��, ��,��^�����������k��g����������_ ��, ��, ��, ��, ��, f�                                                                        ��������-��-������                                                                                                        ������������������                                                                                                        ��
��������������
                                                    ���������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ���������(      0          `	                                                                                                                               p�� p�� o�� n�� m�� l�� k�� j�� j�� j�� j�� j�� j�� j�� j�� j�� i�� U�                         r�� q�� p�� o�� n�� m�� l�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� h�                         s�� r������������������������������������������������������ j�� j�� h�                         t�� t����������������������k������������������������������� j�� j�� h�                         v�� u������������������,]��=��p��������������������������� j�� j�� h�                         w�� v��������������;h��F��T{��@�������������������������� j�� j�� h�                         x�� x����������Eo��A����������O��Hr���������������������� k�� j�� h�                         y�� y������n���@������������������=���������������������� l�� k�� h�                         {�� z������������������������������7e��&X������������������ n�� m�� h�                         }�� |����������������������������������>������������������ o�� n�� h�                         ~�� }����������������������������������]���F�������������� p�� p�� h�                         �� ~��������������������������������������F��a����������� r�� q�� h�                         ��� �������������������������������������������>���������� s�� r�� h�                         ��� �������������������������������������������$V��;h������ t�� t�� h�                         ��� �����������������������������������������������_������� v�� u�� t�                         ��� ������������������������������������������������������� w�� v�� t�                         ��� ������������������������������������������������������� y�� x�� t�                         ��� ���������������@���.���.���.���.���.���.��������������� z�� y�� t�                         ��� ���������������_���c���`���]���Z������}�������� {�� z�� s�                         ��� ��� ��� ��� ������"���"���"���"���!������w�� ��� ��� ��� ��� w�                         �� ��, ��, ��, ��,��g��������@��������o ��/ ��, ��, ��, w�                                                    ���������������                                                                            �������������"                                        ��� �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ��� ��� (      (          �                                                                                                               p�� o�� n�� m�� k�� k�� j�� j�� j�� j�� j�� j�� j�� j�� U�                     r�� q�� p�� o�� n�� m�� k�� j�� j�� j�� j�� j�� j�� j�� h�                     t�� s������������������������������������������ j�� j�� h�                     u�� t��������������l���F���������������������� j�� j�� h�                     w�� v����������{���>��J��T{������������������ j�� j�� h�                     x�� x����������=����������=������������������ l�� k�� h�                     {�� y������$V�������������>j��-]�������������� m�� l�� h�                     |�� {��������������������������>�������������� o�� n�� h�                     ~�� }��������������������������g���J���������� q�� p�� h�                     ��� ������������������������������I��m������� s�� q�� h�                     ��� �����������������������������������@������ t�� s�� h�                     ��� �����������������������������������[������� v�� u�� t�                     ��� ������������������������������������������� x�� v�� t�                     ��� ������������������������������������������� y�� x�� t�                     ��� �����������@���.���.���.���.���.����������� {�� z�� p�                     ��� ������������_���b���^���[������������ ��� ��� y�                     �� ��, ��, ��,���"���!���!���!��������8 ��, ��, y�                                            ������������                                                                ��S��������f                                ��� � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � 0 � p �� �� (                 @                                                                                           p�� o�� n�� l�� k�� j�� j�� j�� j�� j�� j�� f�
                 r�������������������������������������� j�� h�                 u�������������������������������������� j�� h�                 w��������������P��F������������������ j�� h�                 y����������&X��e���Px��]��������������� k�� h�                 {����������[�����������D�������������� m�� h�                 }����������������������w���7e���������� o�� h�                 ��������������������������O���������� q�� h�                 �������������������������������O������ s�� h�                 �������������������������������Ir������ u�� t�                 ��������������������������������������� w�� t�                 �����������@���7���6���5���/����������� y�� t�                 ������������C���A���?��� ��������� �� z�                 |�! ��, ��,��Y�����l�����` ��. ��, |�!                                    ���������                            ��  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  
KeyPreview	PositionpoOwnerFormCenterOnAfterMonitorDpiChangedFormAfterMonitorDpiChangedOnShowFormShow
TextHeight TPanelPanelLeft2Top Width� Height�AlignalRight
BevelOuterbvNoneConstraints.MinHeight^TabOrder
DesignSize� �  TButtonOkButtonLeftTopWidthwHeightAnchorsakLeftakTopakRight CaptionOKDefault	ModalResultTabOrder OnClickOkButtonClickOnDropDownClickOkButtonDropDownClick  TButtonCancelButtonLeftTop'WidthwHeightAnchorsakLeftakTopakRight Cancel	CaptionAvbrytModalResultTabOrder  TButtonCheckAllButtonLeftTop� WidthwHeightActionCheckAllActionAnchorsakLeftakTopakRight TabOrder  TButtonUncheckAllButtonLeftTop� WidthwHeightActionUncheckAllActionAnchorsakLeftakTopakRight TabOrder  TButtonCheckButtonLeftTopuWidthwHeightActionCheckActionAnchorsakLeftakTopakRight TabOrder  TButtonUncheckButtonLeftTop� WidthwHeightActionUncheckActionAnchorsakLeftakTopakRight TabOrder  TButton
HelpButtonLeftTopFWidthwHeightAnchorsakLeftakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TButtonCustomCommandsButton2LeftTop?WidthwHeightActionCustomCommandsActionAnchorsakLeftakTopakRight Caption
Ko&mmandonTabOrder	  TButtonReverseButtonLeftTopWidthwHeightActionReverseActionAnchorsakLeftakTopakRight TabOrder  TButtonToolsMenuButtonLeftTopnWidthwHeightAnchorsakLeftakTopakRight Caption&VerktygTabOrder
OnClickToolsMenuButtonClick  TButton
MoveButtonLeftTop WidthwHeightAction
MoveActionAnchorsakLeftakTopakRight TabOrder   TIEListViewListViewLeft Top Width2Height�
OnRecreateListViewRecreateAlignalClient
Checkboxes	Constraints.MinWidth� DoubleBuffered	FullDrag	HideSelectionReadOnly		RowSelect	ParentDoubleBufferedParentShowHint	PopupMenuListViewPopupMenuShowHint	TabOrder OnChangeListViewChange
OnChangingListViewChangingOnClickListViewClick
NortonLikenlOffColumnsCaptionNamnMaxWidth�MinWidth CaptionLokal katalogMaxWidth�MinWidthWidthd 	AlignmenttaRightJustifyCaptionStorlekMaxWidth�MinWidthWidthF Caption   ÄndradMaxWidth�MinWidthWidthP MaxWidthMinWidthWidth Caption   FjärrkatalogMaxWidth�MinWidthWidthd 	AlignmenttaRightJustifyCaptionStorlekMaxWidth�MinWidthWidthF Caption   ÄndradMaxWidth�MinWidthWidthP  	ViewStylevsReportOnAdvancedCustomDrawSubItem!ListViewAdvancedCustomDrawSubItem	OnCompareListViewCompareOnContextPopupListViewContextPopupOnSelectItemListViewSelectItemOnSecondaryColumnHeaderListViewSecondaryColumnHeader  
TStatusBar	StatusBarLeft Top�Width�HeightHint9   Klicka för att markera alla åtgärder av den här typenPanelsStylepsOwnerDrawText'   Fullständiga synkroniseringsåtgärderWidth_ StylepsOwnerDrawTextNya lokala filerWidth_ StylepsOwnerDrawText   Nya fjärrfilerWidth_ StylepsOwnerDrawTextUppdaterade lokala filerWidth_ StylepsOwnerDrawText   Uppdaterade fjärrfilerWidth_ StylepsOwnerDrawText   Gamla fjärrfilerWidth_ StylepsOwnerDrawTextGamla lokala filerWidth_ Width2  ParentShowHintShowHint	OnMouseDownStatusBarMouseDownOnDrawPanelStatusBarDrawPanelOnResizeStatusBarResize  TPngImageListActionImages	PngImages
BackgroundclWindowName'Total actions counter on sync checklistPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:51+01:00" xmp:MetadataDate="2022-09-01T11:02:51+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:47e94351-a6d1-0049-8587-acbdc6ac7222" xmpMM:DocumentID="adobe:docid:photoshop:8467c3b1-44c7-774c-9258-74380922199f" xmpMM:OriginalDocumentID="xmp.did:58152de4-4f2f-b54d-b050-26bde3c0f9c4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:58152de4-4f2f-b54d-b050-26bde3c0f9c4" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:47e94351-a6d1-0049-8587-acbdc6ac7222" stEvt:when="2022-09-01T11:02:51+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  �IDATxڝ�_HSQ���*����*����0�'2�����՛�Pk�J��oR���C``�d�m1-��� !
��i�ڟ����y�+�������w����9��z����.�\�zW��0Dv��୛�X�q�~y_Y��GV��AxYi��u�^[#n��H0;L	�$}|�n
Kj�6��X	�?5�HK7YE��a^4\ץf��z8����/p�{��~���
k�M��>��X
�cF�� q�;?�8t;���̘
� 3�ć����	,�����s��@"&����%n��8�@�t-JO� �w�[BR1�\#n��+c#��������y�8Ą	𺇸�WEx|�����G�XG&P|�9��Ӌ�����J�ҧ"��Bg����Z( �PA�w<����[p�W���d~!�}A��E��O�VY����L���[������c���}ә�����׷~Hy�'N��i(է"CϿKƈ����8�	��XB+$�"WW�    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:54+01:00" xmp:MetadataDate="2022-09-01T11:02:54+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:a531e4a3-3e94-7044-8248-c5109dce3d50" xmpMM:DocumentID="adobe:docid:photoshop:5ed61c57-dde9-3142-9e44-3c21d266d6a5" xmpMM:OriginalDocumentID="xmp.did:d99e8793-8092-5a44-b637-16371014aa2a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d99e8793-8092-5a44-b637-16371014aa2a" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:a531e4a3-3e94-7044-8248-c5109dce3d50" stEvt:when="2022-09-01T11:02:54+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>R��   �IDATx�c���?%�q@�����>������y����߿����|�7 "���? ��:|�*s��?��1Pn��/��6�2|c�9����.���E�@�����p����xƨ}��Wz|�.v � ���#v!��*�OX�"�! s�~�\�:��с�h���/��cLZ�����w��o�S6�E����7  �g����L�    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:57+01:00" xmp:MetadataDate="2022-09-01T11:02:57+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f42fbb72-a7b3-6c40-a941-b37179109e79" xmpMM:DocumentID="adobe:docid:photoshop:d0604d78-47ae-2942-a011-b611af95bfee" xmpMM:OriginalDocumentID="xmp.did:894a1a4c-b18d-c44c-9f30-83fe31bf3c38"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:894a1a4c-b18d-c44c-9f30-83fe31bf3c38" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f42fbb72-a7b3-6c40-a941-b37179109e79" stEvt:when="2022-09-01T11:02:57+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>D�3�   �IDATx�c���?%�q�.{�C����p��<��:���8�����b���D��[���y##�'#H�����_�G��3]fd*b
21\���/�c�.�P&&�Y@� H3� ��W�|���S�@C��1�o�	e`a�4P �����W~|���
T����WL1��X� mw�y��6V&��0CA����)���;����8	(qo��g��E&�ҕ蓐�� Ȅi�UUvD    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:01+01:00" xmp:MetadataDate="2022-09-01T11:03:01+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ec66effc-45b6-7040-8709-7f0e8e4388fd" xmpMM:DocumentID="adobe:docid:photoshop:072a6ef4-2973-824a-a7bb-58f69dc582d4" xmpMM:OriginalDocumentID="xmp.did:fc555fcc-ee49-124b-aea0-99e4d6ef7c7f"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:fc555fcc-ee49-124b-aea0-99e4d6ef7c7f" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ec66effc-45b6-7040-8709-7f0e8e4388fd" stEvt:when="2022-09-01T11:03:01+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�X�0   �IDATx�c���?%�q@��'a�~��������x"����/��������v�OB���������`���#V�G�� @�߿s߽��gr���C�� E0ʻp��	 �� 3h����3���������.��u��f����Mf�������*vσn Pn��?�0|!:�r�g���ş�����E"��vd[�������8�)q�  ���7�e�    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:05+01:00" xmp:MetadataDate="2022-09-01T11:03:05+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:90325f3a-6b16-a048-8c6e-51cf34e29d43" xmpMM:DocumentID="adobe:docid:photoshop:96bc9090-deaf-9b43-94f8-f83e65f4f27f" xmpMM:OriginalDocumentID="xmp.did:9cc5bf16-41fd-4844-83d8-6e3cbd770e47"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:9cc5bf16-41fd-4844-83d8-6e3cbd770e47" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:90325f3a-6b16-a048-8c6e-51cf34e29d43" stEvt:when="2022-09-01T11:03:05+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��H   �IDATx�ݒ�A�g玓C�]Is�V):A�W����B�/��JT���hw���H$l2���~3;����%� �(ڹ����m�6�����2`�L{²fL�`"`�2QHB�!+sV&$f�&��\W�ژ���:�Lf݀�&�"(�Dډib��t!pn C��Hp�F�5s�M<�N͵�n��C��� ��J�$�vL��j��x��;M��R�:8�W���G�}�~R��
��A    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:11+01:00" xmp:MetadataDate="2022-09-01T11:03:11+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8695f242-2b65-2240-9085-8a3d5c3b269e" xmpMM:DocumentID="adobe:docid:photoshop:96151f7f-c345-e242-be87-01ac864bf8ca" xmpMM:OriginalDocumentID="xmp.did:98a7e7ee-2b00-5347-966c-576201d69420"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:98a7e7ee-2b00-5347-966c-576201d69420" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8695f242-2b65-2240-9085-8a3d5c3b269e" stEvt:when="2022-09-01T11:03:11+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>@Yk  ~IDATxڥ�=K�@��Kb� �"Zď�~D��ͥ]t�{��\�C���Gd��"�`t�"�����K��6ѡ!p���CDXf1-�o{N��H�Zի~���X���_Q�<�~�F�v��ӿJ�*ND�z��6��Y�vnBaË�}*�CT!�rA2��@�n�=0�ζ88��&�Dm,)�k��as�^Z��"	���I,����j
����F!HB���Iʖ����3���q�fN��(����:2@<xZ�Rލ�K��u� �n#��I�'�_�"8���d��8�י�ۑ�$�^c���m$���Kl3� ��C��kcӧ3�2x*q�%�@�ۿ��F��tͫ8nӨ5��ɱ˩�T��1{Lˬ��y�ήO�    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:08+01:00" xmp:MetadataDate="2022-09-01T11:03:08+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f0f22f02-53ea-d145-b8d1-3eb048630a1c" xmpMM:DocumentID="adobe:docid:photoshop:b996e4e5-69df-1e4f-9c5d-d89b233a8f06" xmpMM:OriginalDocumentID="xmp.did:38bc3802-b617-5547-a3cb-91930445c2c8"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:38bc3802-b617-5547-a3cb-91930445c2c8" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f0f22f02-53ea-d145-b8d1-3eb048630a1c" stEvt:when="2022-09-01T11:03:08+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�pyZ  ~IDATxڥ�=K�@��Kb� �"Zď�~D��ͥ]t�{��\�C���Gd��"�`t�"�����K��6ѡ!p���CDXf1-�o{N��H�Zի~���X���_Q�<�~�F�v��ӿJ�*ND�z��6��Y�vnBaË�}*�CT!�rA2��@�n�=0�ζ88��&�Dm,)�k��as�^Z��"	���I,����j
����F!HB���Iʖ����3���q�fN��(����:2@<xZ�Rލ�K��u� �n#��I�'�_�"8���d��8�י�ۑ�$�^c���m$���Kl3� ��C��kcӧ3�2x*q�%�@�ۿ��F��tͫ8nӨ5��ɱ˩�T��1{Lˬ��y�ήO�    IEND�B`�  Left0Top�  
TPopupMenuListViewPopupMenuLeft�Top� 	TMenuItem	CheckItemActionCheckAction  	TMenuItemUncheckItemActionUncheckAction  	TMenuItemN3Caption-  	TMenuItemCheckAllFilesinThisDirectory1ActionCheckDirectoryAction  	TMenuItem!UncheckAllActionsinThisDirectory1ActionUncheckDirectoryAction  	TMenuItemN1Caption-  	TMenuItemReverseItemActionReverseAction  	TMenuItemMoveItemAction
MoveAction  	TMenuItem
Calculate1ActionCalculateSizeAction 	TMenuItem
Calculate3ActionCalculateSizeAction  	TMenuItemCalculateAll1ActionCalculateSizeAllAction   	TMenuItem ActionCustomCommandsAction 	TMenuItem    	TMenuItemBrowseLocalDirectory2ActionBrowseLocalAction  	TMenuItemBrowseLocalDirectory1ActionBrowseRemoteAction  	TMenuItemN2Caption-  	TMenuItemSelectAllItemActionSelectAllAction   TTimerUpdateTimerEnabledIntervaldOnTimerUpdateTimerTimerLeftPTop�  TActionList
ActionListLeft�Top� TActionUncheckActionCaption	Avmarkera	OnExecuteUncheckActionExecute  TActionCheckActionCaptionMarkera	OnExecuteCheckActionExecute  TActionCheckAllActionCaptionMarkera &alla	OnExecuteCheckAllActionExecute  TActionUncheckAllActionCaptionAvmarkera a&lla	OnExecuteUncheckAllActionExecute  TActionSelectAllActionCaption&Markera allaShortCutA@	OnExecuteSelectAllActionExecute  TActionCustomCommandsActionCaptionEgna ko&mmandon	OnExecuteCustomCommandsActionExecute  TActionReverseActionCaption   &Omvänt	OnExecuteReverseActionExecute  TActionCalculateSizeActionCaption	   B&eräknaShortCut�  	OnExecuteCalculateSizeActionExecute  TActionCalculateSizeAllActionCaption   Beräk&na allaShortCut�  	OnExecuteCalculateSizeAllActionExecute  TAction
MoveActionCaption&FlyttaShortCutu	OnExecuteMoveActionExecute  TActionCheckDirectoryActionCaption(   Markera alla åtgärder i &denna katalog	OnExecuteCheckDirectoryActionExecute  TActionUncheckDirectoryActionCaption*   Avmarkera alla åtgärder i denna &katalog	OnExecuteUncheckDirectoryActionExecute  TActionBrowseLocalActionCaption   Bläddra &lokal katalog	OnExecuteBrowseLocalActionExecute  TActionBrowseRemoteActionCaption   Bläddra &fjärrkatalog	OnExecuteBrowseRemoteActionExecute  TActionFindMoveCandidateActionCaption&Hitta flyttkandidatShortCutu�  	OnExecuteFindMoveCandidateActionExecute   TPngImageListActionImages120HeightWidth	PngImages
BackgroundclWindowName'Total actions counter on sync checklistPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:52+01:00" xmp:MetadataDate="2022-09-01T11:02:52+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:acc73d43-b0ee-a647-a8e2-5103fa7f4789" xmpMM:DocumentID="adobe:docid:photoshop:912058f6-e783-494a-941a-e2b245a6d850" xmpMM:OriginalDocumentID="xmp.did:26f8ffbb-3b7d-c546-9636-f483276b3601"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:26f8ffbb-3b7d-c546-9636-f483276b3601" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:acc73d43-b0ee-a647-a8e2-5103fa7f4789" stEvt:when="2022-09-01T11:02:52+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��  tIDATxڭ�_HSQ������R�ݲD����E��!���7A��z2sM-[��=D�b�d��c6�9�E�Л�i�_�ܚwN��i��^W���w~��9��&0�A�{]�Qdb=��
���FoT"��@��KZ�@���lJ6���3reߧJ3�0L�9�4g��J����	���d���	)�&��e��`�9��k���4��C2��95�KE�����������H΀�A�﯇�.����	�m� C:|�M��4��<�g��K�G ���gv��j��`�V5R����-O�2��U��B��N�w����3���
��
�@�bnU=|�E�A��c�v�.:���V<��G����vH��zup�����ȹ�+Ҳ����8X�w�����c�<�'�X_Z��Fe��E�,��qR���:�ie�[gBht�;������u�o�yj�25�U�����w��i퀘����lhz������ު�m�
�����#O߬���b��-y�Z��|��J���j�N+oc���s����Q� ){�߁���_.��$I�q��;��F�j��{�
n�n[,�/��0�w�`�?�D������    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
5  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:55+01:00" xmp:MetadataDate="2022-09-01T11:02:55+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c01c71c5-ee28-814d-8e0b-49e6901e72e6" xmpMM:DocumentID="adobe:docid:photoshop:29a80341-e359-fd41-b94e-4da9ee7cd13b" xmpMM:OriginalDocumentID="xmp.did:c4668d4b-97a3-a44a-b4e6-f9346d03dbb2"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c4668d4b-97a3-a44a-b4e6-f9346d03dbb2" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c01c71c5-ee28-814d-8e0b-49e6901e72e6" stEvt:when="2022-09-01T11:02:55+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�q�  IDATx���j�@�g_`��z*(�@5Vϥ��>���ZhP�Ҙ��^<l=(&3�ML��49:0,|��ogvGd��(����pew�eV@etr��5"�r��s�}��RǴ�]h���<�&`��,(U���.e���z�3ΑN����	���6D�Q<2Q���/�CyU>�o�>�ʡј�d�f`�8Z�f]�:���X���zpQ�e"��Q鰾�SjӨB~=_t����m����%u}��f\�qR�͋%���?��,�L�����@    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
5  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:58+01:00" xmp:MetadataDate="2022-09-01T11:02:58+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:93fa1bfa-6b2a-2c48-8586-19426b57bbef" xmpMM:DocumentID="adobe:docid:photoshop:ce31a24c-4e79-1645-9087-bfd007e64cd9" xmpMM:OriginalDocumentID="xmp.did:a0ac05ec-a673-114e-812c-2a4078702317"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:a0ac05ec-a673-114e-812c-2a4078702317" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:93fa1bfa-6b2a-2c48-8586-19426b57bbef" stEvt:when="2022-09-01T11:02:58+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>,��  IDATx�c���?5㨁�1���C"z�ߔ���(60���2 Sq��GF�l``�v�a`b�edbd�/�&������̬����1�^b�	l`���L@10Zu9�8���]��L�Ӏ��!R��b`����p�@�p�������0n �@ ^� ��U�2'��p/���Pdbz���ٕ0�a�����q�vq�Hqh``��ed�_c����!;y�X �F~�+O`��g��Z�R�H9  ��}�ۀ5    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
T  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:02+01:00" xmp:MetadataDate="2022-09-01T11:03:02+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ea562693-3c34-8949-8f21-6c68617225b6" xmpMM:DocumentID="adobe:docid:photoshop:0003f9da-fec0-b14d-970c-ad5e9dc438c5" xmpMM:OriginalDocumentID="xmp.did:2cd4ebb7-2f55-2641-a26e-17660ea896ca"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:2cd4ebb7-2f55-2641-a26e-17660ea896ca" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ea562693-3c34-8949-8f21-6c68617225b6" stEvt:when="2022-09-01T11:03:02+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>��Q  1IDATx���J1�'��EE�ժU_���
*�
�"}�}A|�
�)J}[���ǂI33&#�����c2��0Q�YJM�� �R�2}^�CS)=�L���3�o4y�����q�lm@d,�z[k7v+L��H�_*�$��~�dy�V@n�{k�?� �5D������������,�Ur�J���|�	��lh1����Q��/������ ������cgg6��.��+��F��v����ݟc�Έ��g]-7�L<��^�q�c�m4M+��y+���H_�^!�cg�)0�~�3 �]�9    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
Q  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:05+01:00" xmp:MetadataDate="2022-09-01T11:03:05+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:aa86f0e5-db92-1542-96a1-609f2d24a1e6" xmpMM:DocumentID="adobe:docid:photoshop:603e15e3-f570-1d4b-aeef-d79e6b15ad76" xmpMM:OriginalDocumentID="xmp.did:5f01ea2b-54b8-5a44-8d08-6757e5e17b8e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5f01ea2b-54b8-5a44-8d08-6757e5e17b8e" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:aa86f0e5-db92-1542-96a1-609f2d24a1e6" stEvt:when="2022-09-01T11:03:05+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>;��  .IDATx�c���?5㨁�1���C�'+��͟�(6�/���e@9Eŭ��6����)ї�������X�	�_�3𞗀<�?����2����d��o`�������/�����Xa�G��`��G͞���?>p$��T d������_�?HL3�"tq�����c�ڧ ]�2h�u ���_`��=y�.��j��ý|ÍC�@s,�U;���3�% �~�/Vq�H����"��V���_P�	$�HQ��n�`��iPB�*��	s>AV��G�E�l 5���� �k�yA_�    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:12+01:00" xmp:MetadataDate="2022-09-01T11:03:12+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:075abba9-a96a-4b4a-84d7-e7771dfc4b01" xmpMM:DocumentID="adobe:docid:photoshop:b3cc6734-e412-0540-bd92-2c3b0c4d137f" xmpMM:OriginalDocumentID="xmp.did:feb01262-5f56-6c43-897f-eff3086114a5"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:feb01262-5f56-6c43-897f-eff3086114a5" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:075abba9-a96a-4b4a-84d7-e7771dfc4b01" stEvt:when="2022-09-01T11:03:12+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�+B�  �IDATxڵ��J�@ ����P�E)J���|
��-/�Z<��kjU(z�u)�Է�"b���P463Φ�m�
u!��~��nD$:�o�����o"aah�F�3������>*�׉0 ��V�-	!�C{�Q�	�O78w$�� V��� '"ǭ����S�0��ˣ���  �N�����;��am�ŏ����wP�F�:��7�U3L����8,�P���0��XKЫf1&�k
�Hw���R��a�6�<Bn�l���z~n W�3DmM��*��ɋj���6��s���� 
6��5�������s�m�VT(X��|���j&»_;����#5vVQ���� c�10��NG$�T��%^�D�M�Rj0Ǐs�0?.����߾w����� x1���Dn�VG'{$w�̞;�_���������    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:09+01:00" xmp:MetadataDate="2022-09-01T11:03:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:ff6cfd6c-1aeb-1a41-8f72-95ce8c85597d" xmpMM:DocumentID="adobe:docid:photoshop:cb7fee06-5a66-c447-932a-9cee175f7a8f" xmpMM:OriginalDocumentID="xmp.did:7f82082b-4a62-9343-8a33-9bc4f0f4c585"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:7f82082b-4a62-9343-8a33-9bc4f0f4c585" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:ff6cfd6c-1aeb-1a41-8f72-95ce8c85597d" stEvt:when="2022-09-01T11:03:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����  �IDATxڵ��J�@ ����P�E)J���|
��-/�Z<��kjU(z�u)�Է�"b���P463Φ�m�
u!��~��nD$:�o�����o"aah�F�3������>*�׉0 ��V�-	!�C{�Q�	�O78w$�� V��� '"ǭ����S�0��ˣ���  �N�����;��am�ŏ����wP�F�:��7�U3L����8,�P���0��XKЫf1&�k
�Hw���R��a�6�<Bn�l���z~n W�3DmM��*��ɋj���6��s���� 
6��5�������s�m�VT(X��|���j&»_;����#5vVQ���� c�10��NG$�T��%^�D�M�Rj0Ǐs�0?.����߾w����� x1���Dn�VG'{$w�̞;�_���������    IEND�B`�  Left� Top�  TPngImageListActionImages144HeightWidth	PngImages
BackgroundclWindowName'Total actions counter on sync checklistPngImage.Data
<	  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:53+01:00" xmp:MetadataDate="2022-09-01T11:02:53+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d6f0ad3b-b203-5d4b-bc3a-13271097edfd" xmpMM:DocumentID="adobe:docid:photoshop:0d378041-9634-1f42-8154-f49c9a5f1413" xmpMM:OriginalDocumentID="xmp.did:6f91a7fc-3331-0446-b27c-a0fa79c7f10c"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:6f91a7fc-3331-0446-b27c-a0fa79c7f10c" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d6f0ad3b-b203-5d4b-bc3a-13271097edfd" stEvt:when="2022-09-01T11:02:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>|���  IDATxڭ�_HSQ��͹�T��[Z���HK-�җ
2�"�(�'����o)�`�=�BD=Hf�K��T�E�hdn:]�47�{;�,�t�^�\.�����9�1<��o0WahR(|����x2�˱�>I��	�5� lWp�#��|Ā9F���D͉����Qd���N�)�j2K	+�j@�./'�f&�+�q�$��:~Do�||8��a����Z���bt`��T�{�Q2SBV��?����|��� �m�̳K����d�22�]�#I����3x���Kmg�� :���-� oY -eT�ʁ�%��Jv��<�������b��	����SL#/ ��R �@`�b�"��29B���.��i� �n�ו�]�<0��&oe ����X�(� ;# �*�g��H�9��	P�=��u�S�l �ʘq�� �D�߼���m�������<
XL@o)�J�毟0z!
���P������� z�I��-c�~$k�lk�0���f���3�����l{���Bz�,�7�H���^��l�sWr��T$��}�N��,
L�BKutP`%��c���}@p]7<7l��3ᐨ֓vג�=�X(4�@g>��	��p���f$�j�As��`C4l������R�ȣ����C��Ф�â�ߡ�̼���E�8X�|�,�a�" ��A��e�k�t}�v���,
خ��3���Bh�dޓf�b@����qMy̳.�'��e5�W�{�Z���}���ˣ��?R    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
r  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:56+01:00" xmp:MetadataDate="2022-09-01T11:02:56+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:d243d29b-864b-294d-a152-e5e98841ee24" xmpMM:DocumentID="adobe:docid:photoshop:075b2236-2af6-0f45-a415-703aa33ba41f" xmpMM:OriginalDocumentID="xmp.did:d064948d-bd00-c347-b222-0e0345e51d57"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d064948d-bd00-c347-b222-0e0345e51d57" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:d243d29b-864b-294d-a152-e5e98841ee24" stEvt:when="2022-09-01T11:02:56+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  OIDATx�c���?-�#�J�;η���OY�}���~` �����߈�v_/Q݂أ`��������/3Q,�� ������������#��c������0�_�����^���] �6B/s�@H>�0�P����;b���S�ч�.��Pb�p�@P� T�ɒ ��/ ��1j?Ȇ�t�@H>� � ��_@�W3F�*��n;�*/��� ����;l�0�"vA]�.	0�G�C�����?�}N����*�4r,�������j�/S��"v-`��ϟak=i��"v�.���s��0�/��Ai:j��[  COJ$��f    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:59+01:00" xmp:MetadataDate="2022-09-01T11:02:59+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:f1002cdf-fd53-0f4b-95dc-ab6c52dfe0f7" xmpMM:DocumentID="adobe:docid:photoshop:8817b227-0de1-f443-97b3-3f3fecac8789" xmpMM:OriginalDocumentID="xmp.did:e72a4056-1ad1-684d-9f4e-55c729afc832"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:e72a4056-1ad1-684d-9f4e-55c729afc832" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:f1002cdf-fd53-0f4b-95dc-ab6c52dfe0f7" stEvt:when="2022-09-01T11:02:59+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  hIDATx�c���?-�#�\���8��[�׹����Zu�C���m#�ÿ�⋭����1�x��� eA�T��a?�_7P $
6L�[}��%�#gb���!.y���x�YV]��j8��o��׻y���%#� &L�������8(��n8���bA�n�0�0��}�/� (1(��n8���b@�ޗ@����� j���/��-<���+�\=��0�0B�@r!Ԑ��#"y>����o�����7� `���SR8���_#����	fbb���)��b U3Z�NE`F[�5����-L���~2�o�������n �U��@V3	    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:03+01:00" xmp:MetadataDate="2022-09-01T11:03:03+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c10af81e-07f1-6549-a519-c43636a259bf" xmpMM:DocumentID="adobe:docid:photoshop:8ebbe314-6816-1c44-bd52-9408929eafe7" xmpMM:OriginalDocumentID="xmp.did:6f85f4d1-1437-784e-a84f-a12720cee115"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:6f85f4d1-1437-784e-a84f-a12720cee115" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c10af81e-07f1-6549-a519-c43636a259bf" stEvt:when="2022-09-01T11:03:03+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�T~h  nIDATx�c���?-�#�Jx&����Y&���Ă'�b���������M�/Q݂����P���������7~��b��0q�<P��� ��3(l������@a���k�������؂�A"�a��P��l !��B� B� ��1��P����C?A���3 ���;� ����b ���������_�xߛŅP���_`�?��; a�����s�g���� $ߋ�����=���_���ߧ�8s��
`������zh0������_)�>P%��u�Y��R�}��P5�q�������߿��i�E��vˑm����r�0|�&?J�Q� �T�4����    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
�  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:06+01:00" xmp:MetadataDate="2022-09-01T11:03:06+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:38844115-f9d9-2c4b-8186-2091eac66d2b" xmpMM:DocumentID="adobe:docid:photoshop:6ffaf430-97df-454c-9e77-d60294a45118" xmpMM:OriginalDocumentID="xmp.did:8c088b8e-f078-f64f-8dfd-69fdf7559e21"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:8c088b8e-f078-f64f-8dfd-69fdf7559e21" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:38844115-f9d9-2c4b-8186-2091eac66d2b" stEvt:when="2022-09-01T11:03:06+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���  �IDATx�픿K�P�/���ml1��R("ԭ� ((,�]�7����8�s�࢓�� ER:���i�����t�{^�}���ܽ<	a�!M � �%<��?�9mT�Y���1R��
.*�?���ŵ�m�22��^$�Ժ(��*����p� O�s�! GC ޏ�2"�G�	����L|��. ���}r��	rv� ��{����\�s�:+g5Q��.���p��#��cl]�aZ�J�2��*{5LQ��.w���+�O��S�PL��� \-�7�CuѢEQ|9rL8��&���v�*���P�7�;�� �c��v[�l���x�Ǵ���){C�3n���h�IX�J�^�c�a_S�rL��?������N ��4ҭ�t��    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
b  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:13+01:00" xmp:MetadataDate="2022-09-01T11:03:13+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:21b8a380-0124-7a40-9ac1-7dd087f2867d" xmpMM:DocumentID="adobe:docid:photoshop:2ebb6369-6404-f545-9ee2-d6da2398c37a" xmpMM:OriginalDocumentID="xmp.did:bfcda6fb-158b-ee4a-bb9d-82e4253090d2"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:bfcda6fb-158b-ee4a-bb9d-82e4253090d2" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:21b8a380-0124-7a40-9ac1-7dd087f2867d" stEvt:when="2022-09-01T11:03:13+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>e���  ?IDATxڽ��n�@�g�4���5=�V	��|@=aY�U�3�7��"������Gh8s�*��N�m��ìc�6n�(�e���3�k��0͇�7c~�Y� �{��W+���ޮ� ��w���V�M�tޮi�4����N�5꒒�`� y����C����)�h�:u�n�d�8��ヽ3#/x�����xb49��#%7����9��~��P��T�J�a�
-�����<�~�P!H�*e�b4��%&����]�7���G�6J� �J&�f��t��&@�����
RI��k(Qa�!���a��8z.%HS�h��+���K2H�m��$x4|rA�s��$Pla���c��@���:d�q�Dq�E��������#������DE�u]�����1���r�t<���zW���SM��d��*�DQ�-��[x���R���+��e'�J��J�
j	�V�����G��߶k�	�!�J�s�I)HWB��>��s��%af��eYxVR)U��j ���pD�>_4fgػ���B���V�yr�?��z�.�jȌ�ENA    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
b  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:09+01:00" xmp:MetadataDate="2022-09-01T11:03:09+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:e4b15b72-9075-db43-a479-979fb0c01f8c" xmpMM:DocumentID="adobe:docid:photoshop:72796009-e0de-d74d-a1a2-3711379443d9" xmpMM:OriginalDocumentID="xmp.did:fead0be8-1316-7046-b1c1-04c7909d5ffd"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:fead0be8-1316-7046-b1c1-04c7909d5ffd" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:e4b15b72-9075-db43-a479-979fb0c01f8c" stEvt:when="2022-09-01T11:03:09+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>w��  ?IDATxڽ��n�@�g�4���5=�V	��|@=aY�U�3�7��"������Gh8s�*��N�m��ìc�6n�(�e���3�k��0͇�7c~�Y� �{��W+���ޮ� ��w���V�M�tޮi�4����N�5꒒�`� y����C����)�h�:u�n�d�8��ヽ3#/x�����xb49��#%7����9��~��P��T�J�a�
-�����<�~�P!H�*e�b4��%&����]�7���G�6J� �J&�f��t��&@�����
RI��k(Qa�!���a��8z.%HS�h��+���K2H�m��$x4|rA�s��$Pla���c��@���:d�q�Dq�E��������#������DE�u]�����1���r�t<���zW���SM��d��*�DQ�-��[x���R���+��e'�J��J�
j	�V�����G��߶k�	�!�J�s�I)HWB��>��s��%af��eYxVR)U��j ���pD�>_4fgػ���B���V�yr�?��z�.�jȌ�ENA    IEND�B`�  Left� Top�  TPngImageListActionImages192Height Width 	PngImages
BackgroundclWindowName'Total actions counter on sync checklistPngImage.Data
�	  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:53+01:00" xmp:MetadataDate="2022-09-01T11:02:53+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:1c48e6a1-7b46-c845-88b7-429fe6da7692" xmpMM:DocumentID="adobe:docid:photoshop:7bbddab3-0cdd-6842-8a9d-695d3d1e8d59" xmpMM:OriginalDocumentID="xmp.did:026e59c7-eb06-614a-b605-1b6d07275072"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:026e59c7-eb06-614a-b605-1b6d07275072" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:1c48e6a1-7b46-c845-88b7-429fe6da7692" stEvt:when="2022-09-01T11:02:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�o(  �IDATx���YLA��R)x!�����x�CPD���4�x'(P�r#P0�xĨ��/��QNi�>�@4F��ҢH@-t�݆�Z���K63����d:�-ò,F�00��!�?]�if�[�K��$s�L~�%��ji>�Ef<9
�BT	�����q��\/ab��a�v�`���+\�Ķ�,�l}f�O_���q`S�4����_�XP�2߹b�輧�4�P�Q�u:��Iah���y��=�Rt�����K��ԶU��
..���Kdd��� ����Z��l�#(��g����0�jԋ_B��,ԟd���\+�[*a/�B�	`S�8|�����Q�F !
J@sx'Xx�J ��)�ΐ�O�� �v �p�+�D�0<J!��J@S6I�N��T���,H�)!�X�:9���<�"i�dz�P����ar�n��]r��b�Q?G	h�$i?9=�Cq}M�p/i���!W�D [�S�d���:���P����<L��1�	`k!%�!��צR �Ϊc�����-�sWdh�J �m(�i�4������0+�&��l�V)#��E��ǩ�>C`�{��O�x.�1j1���LE٘�����"%�Q
dj���c!)����V��!Ƿ;Ep+n��ǘ����K��:9fi���:&C]_ �X�	n�~��w�t`v�����SK �)���![��W��Ң:�\��Y!|��c�L�jP~J��*n�]W(5I�����GM4��Q�����gJ�~�*�bĆ:5�:� �r�O���+�N@��񼥘}�9��gU	�;��*�ջ�݂�"/�� �2ؔg�ϱE�������X�B2�l�>�&��O�@Ԁ�������'V="���
�/�~��u���Uy    IEND�B`� 
BackgroundclWindowNameNew local files indicatorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:02:57+01:00" xmp:MetadataDate="2022-09-01T11:02:57+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c8de9864-1251-0143-973a-616bfca2eba6" xmpMM:DocumentID="adobe:docid:photoshop:ac72b163-c17e-1d43-bc18-116260247203" xmpMM:OriginalDocumentID="xmp.did:52700f95-ad6f-8944-9f16-d09fb35a0543"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:52700f95-ad6f-8944-9f16-d09fb35a0543" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c8de9864-1251-0143-973a-616bfca2eba6" stEvt:when="2022-09-01T11:02:57+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>x���  �IDATx���N�@�O�����AL\�E�M����ְr�x)5Wމ(����L�A+���qz����5!�p&��i���o�LgD�Q�p �m�|��ڭ�J>�Y@EҒ�H��m%[�:T�DYB0g����vƕR_�dU2��Y�=ϻ�7ү.q���v!ۄ@J*�= ��m��^�4����т��*�䒒�4Eb ��ېEy�i���$ڙ���e��Ey����o��Y;?e�Ugi��MU���d�X����C��_]��S�h[YA��M|}_b�vʼb!l��݈��k*�(�j�,��)�^�7�Ja�0���A�F����ʖcF�{��3���^�k���r�/H��z��0�be��{M%�t0��F4h�ȅhnŘy�(����⹳����'!���ȏc�8�����A�    IEND�B`� 
BackgroundclWindowNameNew remote files indicatorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03+01:00" xmp:MetadataDate="2022-09-01T11:03+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:bbfe10dd-8fad-b64e-a848-b386a98970cf" xmpMM:DocumentID="adobe:docid:photoshop:04eaf632-f16f-854d-ab5b-981d9179d6f6" xmpMM:OriginalDocumentID="xmp.did:99de3a80-3222-6f41-8d68-c04d71633f38"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:99de3a80-3222-6f41-8d68-c04d71633f38" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:bbfe10dd-8fad-b64e-a848-b386a98970cf" stEvt:when="2022-09-01T11:03+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�'��  �IDATx��MKQ�Ϲ����h���6A���PDP�Z�h-�
B��~���j#�&���{�zgD�Q]4�s�yy�9����D�� , �0+T>s6���p� �2H�L�3��,g6�c�� JE^�!<����G .�>� ���{I\��[ ��^1>�3"5���ߜ� 	,�/��-�aZ��� �)�Ͼ�dd�em��Z �k�{�U�tT�}$�:�%�O?=dd��܆9��=���x�_.�o��:�-��Ucc=� ]���>h�@_u{+
;�8Rƽ�3�k� Rr-�%����꺰��{����麆PY�Cx�S�l$�8��۸Ő9��g��,���-��2VJ���aV��P9yqA�{��Hg<�|'A�Y�〘�b���8z���О.�jC���� ,����7�g�    IEND�B`� 
BackgroundclWindowNameModified local files indicatorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:04+01:00" xmp:MetadataDate="2022-09-01T11:03:04+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:550cf6ba-f3ab-5f45-84b0-c9c3640528c8" xmpMM:DocumentID="adobe:docid:photoshop:21ddce43-e13b-a248-b1e9-3cc322f12ebc" xmpMM:OriginalDocumentID="xmp.did:c9f70539-0051-1848-a129-a3c8ec5ed16e"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:c9f70539-0051-1848-a129-a3c8ec5ed16e" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:550cf6ba-f3ab-5f45-84b0-c9c3640528c8" stEvt:when="2022-09-01T11:03:04+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>���g  �IDATx��KKQ��lBJzP�"���5��AQDQ}�H�6�.(܆��-��QB���u��,Swf�h:��ә;3���.���������=�� ie�, �� m�Zw������y&����<i?�~���Dl.�J?�i���q�������(��������4�K,�� �PJ�?.d%̦k Hld�����I��R/(�5���i��9�~�� #C�}�2W66��/��R�J mJ ��Q��@|�@5�2�dr�*(��A�R	ym���+JE/�2�	ՆLPN4v+0c����.З��
ecZ��b3v02��!���U�֌^Y?�H6���<O��"�D���Ƈ%flV�����'��ܔ��at����Pk��Y]l���Ɲ�p��m�胈UJ�h���;��A�h��������MR��G�팓�-g����Z~[ ���~ N-�Kz��    IEND�B`� 
BackgroundclWindowNameModified remote files indicatorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:07+01:00" xmp:MetadataDate="2022-09-01T11:03:07+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:caf4a560-1c86-374b-805b-f091f8665524" xmpMM:DocumentID="adobe:docid:photoshop:d3a46e3d-eb2b-ba4c-a5b4-bcf2299eb5d0" xmpMM:OriginalDocumentID="xmp.did:3f67468b-b1c9-754f-a6b3-09d3da8cf673"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:3f67468b-b1c9-754f-a6b3-09d3da8cf673" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:caf4a560-1c86-374b-805b-f091f8665524" stEvt:when="2022-09-01T11:03:07+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>+���  �IDATx�c���?�@�Q�:`�� V�7NYVv���?���Xx�K��3�����Kq�'�M�y���gd��&pD�Kq�g�;�/�s��xpb�����X��p����Aš��� j�|�-�R���D�d���r!��ȎP����q��l���B��:���q�1�g����������Uv�y(���0��ίD�c������+����`�5r���6������P�PZv��ԁ����
,��|_�������������j ����Xu�(���m���8�Ȃ��ȎP;����l�,R?�(u�0ƅ#�����cq��n\�!��c@O� �~�/Q�gCFF��d<��h�q� '.ta�Xux��,��p� B7��2����"e�TTX��������kV�,L̓Վ�����:u��F0�  �H8�U��    IEND�B`� 
BackgroundclWindowNameObsolete local files indicatorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:13+01:00" xmp:MetadataDate="2022-09-01T11:03:13+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:2bf23562-8965-264c-be80-129617eea08b" xmpMM:DocumentID="adobe:docid:photoshop:e0fceecd-dd84-1f4b-a606-b89566ebf534" xmpMM:OriginalDocumentID="xmp.did:a2f57263-e0e4-b64e-9abd-15819a0af257"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:a2f57263-e0e4-b64e-9abd-15819a0af257" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:2bf23562-8965-264c-be80-129617eea08b" stEvt:when="2022-09-01T11:03:13+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>v��c  �IDATx���jA�g�-���Ji/�xc�D��"ap���'�"� �b	����BR�U�S% ����3�394�=Ez�!��&����03�~~ �.�9����K�c�6_R_<:�<�n��`��r���x ���M/|��dU�}b�[%V@�魬�ӗ��'���$,� ,�W���H��7��Ü�"�`�6*]��q/�D7�<@�L���Mtܒ�DT��_�?��%���#�N�_�M h	��P�&��o{����0����0㓜�C	`\Kh=Eb��Dxb#AyС4���	'W�zY��ĵ��&�H艙�p'��4��Zb�$8V!)�E��C��Tx&��K�R0�A�;��PQI�,`BM?��)Ф�\V���� �@w��K�T����(o�� �����\�]�����H<�\n-%�g�1�$h���>��S���M�կ�,lQ�5��$��$p3�I�"a�C���c�q#�R�n��>���$�l#���/pw�I#�f�ޒ(H�,8�m�>"I��ߎ���ĥB�X٭<��pg��FH�������!�nƻ�9ġ��~�pn�Y�ed>,�t��ޒ8D��x�sP��h���@}�Xn�[�#Rp���w<�l:��9�_/���x{~d��Ʈ�+R`?Ɓ�?M�X�h\�}    IEND�B`� 
BackgroundclWindowNameObsolete remote files indicatorPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:24+01:00" xmp:ModifyDate="2022-09-01T11:03:10+01:00" xmp:MetadataDate="2022-09-01T11:03:10+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:7e7aa62a-17af-854d-8f4e-248cb8c303bf" xmpMM:DocumentID="adobe:docid:photoshop:382c79bc-8f52-2149-a43e-388a2993b1d0" xmpMM:OriginalDocumentID="xmp.did:16d89670-a484-a44f-b3cf-921e379c685a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:16d89670-a484-a44f-b3cf-921e379c685a" stEvt:when="2022-06-27T15:59:24+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:7e7aa62a-17af-854d-8f4e-248cb8c303bf" stEvt:when="2022-09-01T11:03:10+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�A�_  �IDATx��Mk�@�ߙ� ,(�Xq[7R\/ڃ��AAJ�P�`@Bi�'���H@
�eQDP�UD<� ���*~���[3��L2ُn�l�s�d��<y?ff"�Av(�-�?oݭL�n���Ξ�`�|��{����;[���@딽�d�o�5���Y�V��p�� �ӗ�#�O�$B82NX�-�?������o��A�F�+<!��3�D?\����J����4��I���.W_�
�$�������O'���M�i	T���&ʏ>;���� �����c�3	LI(5Ebi�Dxb-AyP��ϩtЄ�K_�4�����AM��P���Ɨ}��
V4|h%1Gm���jQ˿NO%��rn���(��2*��t�鑞<�M
�$J@���\�s�h�������@4��$aOv�OAT�Ixw ���t'�"ܜ)����V�$h�����C	����<fBТ��@�h�_����po�E"�E����g���=p���jH��P�6-*#�W0����|3J�HM�����r�$~�o�Y�����X�[���aU_�FH�ٓ��px���L�c�Z�,0��]?m�<��'�H�q�T�OY���t���w�h���/���p�K5��|x(qu����%<��tL�2۹�1Y�2r����F_G
�8�]��S�    IEND�B`�  Left8Top�  
TPopupMenuToolsPopupMenuLeftXTopP 	TMenuItem
Calculate2ActionCalculateSizeAction  	TMenuItemCalculateAll2ActionCalculateSizeAllAction  	TMenuItemN4Caption-  	TMenuItemFindMoveCandidate1ActionFindMoveCandidateAction   
TPopupMenuOkPopupMenuLeft� TopP 	TMenuItem	StartItemCaption&StartDefault	OnClickStartItemClick  	TMenuItemStartQueueItemCaptionStarta i &bakgrundenOnClickStartQueueItemClick     TPF0TSynchronizeDialogSynchronizeDialogLeftoTop� HelpType	htKeywordHelpKeywordui_keepuptodateBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaption"Keep remote directory up to date XClientHeight�ClientWidthColor	clBtnFaceFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style 
KeyPreview	PositionpoOwnerFormCenterOnCloseQueryFormCloseQuery	OnKeyDownFormKeyDownOnShowFormShow
DesignSize� 
TextHeight 	TGroupBoxDirectoriesGroupLeftTopWidth�HeightxAnchorsakLeftakTopakRight Caption	KatalogerTabOrder 
DesignSize�x  TLabelLocalDirectoryLabelLeft1TopWidth� HeightAnchorsakLeftakTopakRight Caption.   Be&vaka förändringar i den lokala katalogen:FocusControlLocalDirectoryEdit  TLabelRemoteDirectoryLabelLeft1TopEWidth:HeightAnchorsakLeftakTopakRight Caption6   ... och inför dessa &automatiskt på fjärrkatalogen:FocusControlRemoteDirectoryEdit  TImageImageLeftTopWidth Height AutoSize	  THistoryComboBoxRemoteDirectoryEditLeft1TopWWidth�HeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrderTextRemoteDirectoryEditOnChangeControlChange  THistoryComboBoxLocalDirectoryEditLeft1Top(WidthfHeightAutoCompleteAnchorsakLeftakTopakRight 	MaxLength�TabOrder TextLocalDirectoryEditOnChangeControlChange  TButtonLocalDirectoryBrowseButtonLeft�Top'WidthPHeightAnchorsakTopakRight Caption   &Bläddra...TabOrderOnClickLocalDirectoryBrowseButtonClick   TButton
StopButtonLeft� TopCWidth^HeightAnchorsakTopakRight Caption&StoppTabOrderOnClickStopButtonClick  TButtonCancelButtonLeft<TopCWidth^HeightAnchorsakTopakRight Cancel	Caption   StängModalResultTabOrder  	TGroupBoxOptionsGroupLeftTop� Width�HeightvAnchorsakLeftakTopakRight Caption   Alternativ för synkroniseringTabOrder
DesignSize�v  	TCheckBoxSynchronizeDeleteCheckLeft	TopWidth� HeightCaption&Ta bort filerTabOrder OnClickControlChange  	TCheckBoxSaveSettingsCheckLeft	Top[Width� HeightCaption*   Använd &samma inställningar nästa gångTabOrderOnClickControlChange  	TCheckBoxSynchronizeExistingOnlyCheckLeft� TopWidth� HeightAnchorsakLeftakTopakRight CaptionBara &existerande filerTabOrderOnClickControlChange  	TCheckBoxSynchronizeRecursiveCheckLeft	Top-Width� HeightCaption&Uppdatera underkatalogerTabOrderOnClickControlChange  TGrayedCheckBoxSynchronizeSynchronizeCheckLeft� TopFWidth� HeightAllowGrayed	AnchorsakLeftakTopakRight CaptionSynkronisera vid s&tartTabOrderOnClickControlChange  	TCheckBoxSynchronizeSelectedOnlyCheckLeft� Top.Width� HeightCaption&Bara markerade filerTabOrderOnClickControlChange  	TCheckBoxContinueOnErrorCheckLeft	TopDWidth� HeightCaption   Fortsätt vid &felTabOrderOnClickControlChange   TButtonStartButtonLeft� TopCWidth^HeightAnchorsakTopakRight Caption&StartDefault	TabOrderOnClickStartButtonClickOnDropDownClickStartButtonDropDownClick  TButtonMinimizeButtonLeft<TopCWidth^HeightAnchorsakTopakRight Caption	&MinimeraTabOrderOnClickMinimizeButtonClickOnDropDownClickMinimizeButtonDropDownClick  TButtonTransferSettingsButtonLeftTopCWidth� HeightCaption   Över&föringsinställningarTabOrderOnClickTransferSettingsButtonClickOnDropDownClick#TransferSettingsButtonDropDownClick  	TGroupBoxCopyParamGroupLeftTopWidth�Height;AnchorsakLeftakTopakRight Caption   ÖverföringsinställningarTabOrderOnClickCopyParamGroupClickOnContextPopupCopyParamGroupContextPopup
DesignSize�;  TLabelCopyParamLabelLeft	TopWidth�Height#AnchorsakLeftakTopakRightakBottom AutoSizeCaptionCopyParamLabelShowAccelCharWordWrap	OnClickCopyParamGroupClick   TButton
HelpButtonLeft�TopCWidth^HeightAnchorsakTopakRight Caption   &HjälpTabOrderOnClickHelpButtonClick  TPanelLogPanelLeft TopaWidthHeightqAlignalBottom
BevelOuterbvNoneTabOrder	
DesignSizeq  	TListViewLogViewLeftTopWidth�HeightgAnchorsakLeftakTopakRightakBottom ColumnsWidth�	WidthType�  Width�	WidthType�   DoubleBuffered	ReadOnly		RowSelect	ParentDoubleBufferedShowColumnHeadersTabOrder 	ViewStylevsReportOnCustomDrawItemLogViewCustomDrawItem
OnDblClickLogViewDblClick
OnDeletionLogViewDeletion	OnKeyDownLogViewKeyDown   
TPopupMenuMinimizeMenuLeftxTopx 	TMenuItem	Minimize1Caption	&MinimeraDefault	OnClickMinimize1Click  	TMenuItemMinimizetoTray1Caption   Minimera till system&fältetOnClickMinimizetoTray1Click   
TPopupMenu	StartMenuLeft Topx 	TMenuItemStart1Caption&StartDefault	OnClickStartButtonClick  	TMenuItemStartInNewWindowItemCaption   Starta i &nytt fönsterOnClickStartInNewWindowItemClick     TPF0TSynchronizeProgressFormSynchronizeProgressFormLeftOTopBorderIconsbiSystemMenu
biMinimize
biMaximizebiHelp BorderStylebsDialogCaptionSynchronization XClientHeight� ClientWidth�ColorclWindowFont.CharsetDEFAULT_CHARSET
Font.ColorclWindowTextFont.Height�	Font.NameSegoe UI
Font.Style PositionpoOwnerFormCenter
DesignSize��  
TextHeight TLabelTimeLeftLabelLeft� Top2WidthOHeightAutoSizeCaption00:00:00ShowAccelChar  TLabelTimeLeftLabelLabelLeft2Top2Width2HeightCaption	Tid kvar:ShowAccelChar  TLabelLabel1Left2TopWidthHeightCaptionLokal:ShowAccelChar  TLabelLabel2Left2Top Width,HeightCaption   Fjärr:ShowAccelChar  
TPathLabelRemoteDirectoryLabelLeft� Top WidthHeightUnixPath	IndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  
TPathLabelLocalDirectoryLabelLeft� TopWidthHeightIndentHorizontal IndentVertical AlignalNoneAnchorsakLeftakTopakRight AutoSize  TLabelStartTimeLabelLeft� Top2WidthQHeightAutoSizeCaption00:00:00ShowAccelChar  TLabelStartTimeLabelLabelLeft2Top2Width6HeightCaptionStartad:ShowAccelChar  TLabelLabel3Left2TopDWidthIHeightCaption   Förfluten tid:ShowAccelChar  TLabelTimeElapsedLabelLeft� TopDWidthOHeightAutoSizeCaption00:00:00ShowAccelChar  	TPaintBoxAnimationPaintBoxLeftTopWidth Height   TPanelToolbarPanelLeft2TopsWidth� HeightAnchorsakLeftakBottom 
BevelOuterbvNoneParentColor	TabOrder  TTBXDockDockLeft Top Width� Height	AllowDragColorclWindow TTBXToolbarToolbarLeft Top DockModedmCannotFloatOrChangeDocksDockPos�DragHandleStyledhNoneImages	ImageListParentShowHintProcessShortCuts	ShowHint	TabOrder ColorclWindow TTBXItem
CancelItemCaptionAvbryt
ImageIndex ShortCutOnClickCancelItemClick  TTBXItemMinimizeItemCaption	&Minimera
ImageIndexShortCutM�  OnClickMinimizeItemClick     TPanelComponentsPanelLeft Top� Width�HeightBAlignalBottom
BevelEdgesbeTop 	BevelKindbkFlat
BevelOuterbvNoneTabOrder  TProgressBarOperationProgressLeft2TopVWidthmHeightAnchorsakLeftakTopakRight ParentShowHintShowHint	TabOrder  TTimerUpdateTimerEnabledOnTimerUpdateTimerTimerLeft�Top�   TPngImageList	ImageList	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:34+01:00" xmp:MetadataDate="2022-09-01T10:57:34+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:180c2c88-0c60-ab4a-b417-9c9f76a6e069" xmpMM:DocumentID="adobe:docid:photoshop:b1118248-b8f9-3348-b679-1d9529e70ef5" xmpMM:OriginalDocumentID="xmp.did:d542fc81-8626-f34b-9a93-59aa7ca76804"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:d542fc81-8626-f34b-9a93-59aa7ca76804" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:180c2c88-0c60-ab4a-b417-9c9f76a6e069" stEvt:when="2022-09-01T10:57:34+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�sa  ~IDATxڥ�=K�@��Kb� �"Zď�~D��ͥ]t�{��\�C���Gd��"�`t�"�����K��6ѡ!p���CDXf1-�o{N��H�Zի~���X���_Q�<�~�F�v��ӿJ�*ND�z��6��Y�vnBaË�}*�CT!�rA2��@�n�=0�ζ88��&�Dm,)�k��as�^Z��"	���I,����j
����F!HB���Iʖ����3���q�fN��(����:2@<xZ�Rލ�K��u� �n#��I�'�_�"8���d��8�י�ۑ�$�^c���m$���Kl3� ��C��kcӧ3�2x*q�%�@�ۿ��F��tͫ8nӨ5��ɱ˩�T��1{Lˬ��y�ήO�    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
B  �PNG

   IHDR         ��a   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:49+01:00" xmp:MetadataDate="2022-09-01T11:07:49+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:c268d7f3-d2fb-104b-a1d0-bb0a4d3ff770" xmpMM:DocumentID="adobe:docid:photoshop:2f11441a-416e-0c44-a239-1906973e411c" xmpMM:OriginalDocumentID="xmp.did:f4e92379-e79c-1e49-9b59-46651bc855c3"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:f4e92379-e79c-1e49-9b59-46651bc855c3" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:c268d7f3-d2fb-104b-a1d0-bb0a4d3ff770" stEvt:when="2022-09-01T11:07:49+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>����   IDATx�cd�0�0H�O��0�a0j �  O����.    IEND�B`�  Left(Top�   TPngImageListImageList120HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:35+01:00" xmp:MetadataDate="2022-09-01T10:57:35+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:b6b0eab7-5227-3e4f-b344-ce0b9ec729f8" xmpMM:DocumentID="adobe:docid:photoshop:d07e584c-62e9-1746-8485-b3340c627702" xmpMM:OriginalDocumentID="xmp.did:ffde8c28-ede5-584b-82d1-a4005269b900"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:ffde8c28-ede5-584b-82d1-a4005269b900" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:b6b0eab7-5227-3e4f-b344-ce0b9ec729f8" stEvt:when="2022-09-01T10:57:35+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>/��@  �IDATxڵ��J�@ ����P�E)J���|
��-/�Z<��kjU(z�u)�Է�"b���P463Φ�m�
u!��~��nD$:�o�����o"aah�F�3������>*�׉0 ��V�-	!�C{�Q�	�O78w$�� V��� '"ǭ����S�0��ˣ���  �N�����;��am�ŏ����wP�F�:��7�U3L����8,�P���0��XKЫf1&�k
�Hw���R��a�6�<Bn�l���z~n W�3DmM��*��ɋj���6��s���� 
6��5�������s�m�VT(X��|���j&»_;����#5vVQ���� c�10��NG$�T��%^�D�M�Rj0Ǐs�0?.����߾w����� x1���Dn�VG'{$w�̞;�_���������    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
G  �PNG

   IHDR         ��   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:50+01:00" xmp:MetadataDate="2022-09-01T11:07:50+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:861cdb4d-c261-6245-b6c7-bb3f3ad7f4f0" xmpMM:DocumentID="adobe:docid:photoshop:bab765bc-e4a8-264e-bb48-0f973dcd85cb" xmpMM:OriginalDocumentID="xmp.did:852956c0-5101-6e4b-9e6b-f9cf5676a668"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:852956c0-5101-6e4b-9e6b-f9cf5676a668" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:861cdb4d-c261-6245-b6c7-bb3f3ad7f4f0" stEvt:when="2022-09-01T11:07:50+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>I���   $IDATx�cd�2`5p��Aj�J̠��T�򨁣��@ ���H�    IEND�B`�  Left� Top�   TPngImageListImageList144HeightWidth	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
b  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:36+01:00" xmp:MetadataDate="2022-09-01T10:57:36+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:476080b3-62e3-864e-915a-47b66c957534" xmpMM:DocumentID="adobe:docid:photoshop:182e7d80-cad1-214c-a9e1-1b656de377c2" xmpMM:OriginalDocumentID="xmp.did:581990f0-e9f9-2844-b56d-bd917ec672b0"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:581990f0-e9f9-2844-b56d-bd917ec672b0" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:476080b3-62e3-864e-915a-47b66c957534" stEvt:when="2022-09-01T10:57:36+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>dn  ?IDATxڽ��n�@�g�4���5=�V	��|@=aY�U�3�7��"������Gh8s�*��N�m��ìc�6n�(�e���3�k��0͇�7c~�Y� �{��W+���ޮ� ��w���V�M�tޮi�4����N�5꒒�`� y����C����)�h�:u�n�d�8��ヽ3#/x�����xb49��#%7����9��~��P��T�J�a�
-�����<�~�P!H�*e�b4��%&����]�7���G�6J� �J&�f��t��&@�����
RI��k(Qa�!���a��8z.%HS�h��+���K2H�m��$x4|rA�s��$Pla���c��@���:d�q�Dq�E��������#������DE�u]�����1���r�t<���zW���SM��d��*�DQ�-��[x���R���+��e'�J��J�
j	�V�����G��߶k�	�!�J�s�I)HWB��>��s��%af��eYxVR)U��j ���pD�>_4fgػ���B���V�yr�?��z�.�jȌ�ENA    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
K  �PNG

   IHDR         �w=�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:59:53+01:00" xmp:ModifyDate="2022-09-01T11:07:50+01:00" xmp:MetadataDate="2022-09-01T11:07:50+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:375ecdd0-9fca-6e44-8e6f-e5190740fc98" xmpMM:DocumentID="adobe:docid:photoshop:48e9df4f-c528-184d-bb90-8e84a567edf0" xmpMM:OriginalDocumentID="xmp.did:86b9b7b2-08b0-9f4d-ad35-1e46758e57e4"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:86b9b7b2-08b0-9f4d-ad35-1e46758e57e4" stEvt:when="2022-06-27T15:59:53+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:375ecdd0-9fca-6e44-8e6f-e5190740fc98" stEvt:when="2022-09-01T11:07:50+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>� �   (IDATx�cd�1`�`ԂQƂ��4sxZ@U0j��� �uv�&    IEND�B`�  Left� Top�   TPngImageListImageList192Height Width 	PngImages
BackgroundclWindowNameCancel operationPngImage.Data
�  �PNG

   IHDR           szz�   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?> <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="Adobe XMP Core 7.2-c000 79.1b65a79, 2022/06/13-17:46:14        "> <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#"> <rdf:Description rdf:about="" xmlns:xmp="http://ns.adobe.com/xap/1.0/" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:photoshop="http://ns.adobe.com/photoshop/1.0/" xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/" xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#" xmp:CreatorTool="Adobe Photoshop 23.5 (Windows)" xmp:CreateDate="2022-06-27T15:58:37+01:00" xmp:ModifyDate="2022-09-01T10:57:37+01:00" xmp:MetadataDate="2022-09-01T10:57:37+01:00" dc:format="image/png" photoshop:ColorMode="3" xmpMM:InstanceID="xmp.iid:8ac33e32-9f3e-5048-9d4c-3532138eb0f4" xmpMM:DocumentID="adobe:docid:photoshop:e1d2034c-6c54-f14f-926e-04f6d15de903" xmpMM:OriginalDocumentID="xmp.did:5fa8f5a2-8a46-b542-9d43-49f9de86586a"> <xmpMM:History> <rdf:Seq> <rdf:li stEvt:action="created" stEvt:instanceID="xmp.iid:5fa8f5a2-8a46-b542-9d43-49f9de86586a" stEvt:when="2022-06-27T15:58:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)"/> <rdf:li stEvt:action="saved" stEvt:instanceID="xmp.iid:8ac33e32-9f3e-5048-9d4c-3532138eb0f4" stEvt:when="2022-09-01T10:57:37+01:00" stEvt:softwareAgent="Adobe Photoshop 23.5 (Windows)" stEvt:changed="/"/> </rdf:Seq> </xmpMM:History> </rdf:Description> </rdf:RDF> </x:xmpmeta> <?xpacket end="r"?>�Ǩ�  �IDATx���jA�g�-��̖�^h���(� �E(���g��@|�Ȃ�%PD��荨���Z<������ݙ�͞"���$���������0?h����;7K3#����-����~��ژ��ޚX��s����o��B�Y�^��p�(��t��$�)���#�e������)��un���DL]F�>�3ꦓ��h�/�~����S�)U�*�-� ��Xb�H8�c�~��5����&��@)!kb�᎛Nφ�n��ր��1{�"�+	e��H�v�HO,�%(*��*4���77<���X	k"����)g�Q ��Z@I,��*�� %ԢȜ�wW���$��rq��+��&%dT��3�P�_�B�4)<���`a:2��"Й�E�d.Ml��7�hx�;(�����t�˰Kxgw0jQ��^��p{�h3����M�V���ӊ9!�J�\�w����� �w0$�z��(	\�IP$Lw(R�wL>��_���ܣ�>��`��m[TF�/pg�i=�f�ޔ(�Yph��}D�������`�2[y���L?ۏ>�x�.
��.�!����+{�C�;t�4����ƫ�|�/���rxS��'���@ej��[�\�,8��7��l��<�ߗ��0�;1k�v_���������}3W��a�#�M�X��E��    IEND�B`� 
BackgroundclWindowNameMinimizePngImage.Data
   �PNG

   IHDR           szz�   	pHYs  �  ��o�d   1IDATx���1  �0�_4� ��@�:.      ���xX	     �0��!Hz �    IEND�B`�  Left8Top�      <4   V S _ V E R S I O N _ I N F O     ���   W                                     �   S t r i n g F i l e I n f o   v   0 4 1 D f d e 9   >   C o m p a n y N a m e     M a r t i n   P r i k r y l     n #  F i l e D e s c r i p t i o n     S w e d i s h   t r a n s l a t i o n   o f   W i n S C P   ( S V )     *   F i l e V e r s i o n     1 . 8 7     � 0  L e g a l C o p y r i g h t   �   2 0 0 3  2 0 2 5   A n d r e a s   P e t t e r s s o n   o c h   R e n �   F i c h t e r   < 
  O r i g i n a l F i l e n a m e   W i n S C P . s v   4   P r o d u c t V e r s i o n   6 . 5 . 3 . 0   8   W W W     h t t p s : / / w i n s c p . n e t /   (   L a n g N a m e   S w e d i s h   .   P r o d u c t N a m e     W i n S C P     D    V a r F i l e I n f o     $    T r a n s l a t i o n     ��                                                                                                                                                                                                                                                                                                                                                                                                               �  �9�9v:�=�=�=>M>U>�>�>�>�?�?�?  �788(828<8F88$8.888B8L8X8q8�8�8�8�8�8�8
999'919;9V9_9i9s9}9�9:#:(:Y:^:k:~:�:�:�:�:o;�< ==&=�=E>k>�>�>�>�>?/?9?�?�89Q9�9C3W3l3�3�34(4G4W4x4�4�5�5�5"6�6�6�6�6�6�45@5W5d5t5�5�5�5766�677,737:7A7H7�45�5D6c6h6m6r6�6�6�6�6�6�6�6�6 7U7�7�7�7p7�7�7�700000 0&0,02080>0D0J0P0V0\0b0h0n0�0�0O1d1�0�0�0�0�0�0�0�0�0�0�01"1(111?1H1X1j1{1�1�1�1�12#292B2_2l2z2�2�2�2�2�2�2�2"3+3:3    �   �:�;�;P<Z8�8H:�:�;Y<�8�89�:�:�;<0>z>�89�:�:<<�>89:�<!=�?�9:a;9=}=�?:3:;;W;x;'<�<s=�=�=I>�>�?�?04\5G0R0y0�0�0�2�2�2�2�2 3Q3�3�3�3�3�3555 5-5A5E5K5O5w5~5�5%6760[0c0L2Y2p2�2�213\3|3�3
44%4B4K4�566J6G9N938{8�8h:3<I8�8[: 0  �   �:o;w;�;�;<#<�<�<�<�=�;�;�<�=�=�=�=^;�;�;�;�;�;<0<f<:=�=�=�=�=R>^>?m??�>�>  �0�0:0�0�0U1e1 2202�2�2�2�2 3$3(3,3034383<3@3R4�5�5;6�6�6�6�678'8�8�8~9�9�9�9:B:�:�:	;;;�<:):<:M:e:z:�:�:�:�:�:$;;;�<�<�< @  �   ;;/;C;l<q<�<�<==4=9=q=�=�=�=�=�=�=>->�>�?�>�?�?�0�0�061a1f1t1U0e0�0�0�0�0�0	1101T1�1�1�1;2M2363�3�3�34K3z3�3�3�3�344)4S4�4�4�4555-5t5y5�5U6�6�6�67F7T7]7g7m7w7�7�7�9; P  �   v<�<�<�<�<�<A=L=k=�=�=�= >> >%>(?�?�?6?j011�1$1%282�4T5�3�3�3�3�3�3�3X5_53�45H5j5�56v6�7�7�7�7�7�7�7�7&8,8m8:8�8�8�8G9P9�8�8�8�8k9�9;!;};�:�:�:6;P;];e;k;�;�;�<U<`< `  �   c8s8999"9,99&90999M9�9:�>�9�9�9�<�> ?�?�?�9c;h;;�;�;�;�;.<<<A<�<�<=$=)=L=Q=�=�=�=�=�?�?  0050:0d0i0�0�0�1�1=2B2�2�2�2�2�2�2�23 31363b3g3}3�3�3�3�3�3`5x5�5�5�56[6N6W6a6j6n6u6�6�6�6�6�6�6�6�67$757�7�7.868�8�8�8B8R8 p  �   4;�;�;�;�;�; <?<D<�<�<==�=�=�=�=>!>�>�>  �0�0`4|4060;0�0�0.131M1R1j1o12"2A2F2^2c2�2�2*3/3�3�3�4�4!5/545�5�5�5�5�5%6*677_7d7�7�788�8�8�8�8�9�9�9�9::@:E:e:j:�:�:/; �  �   �7�7�7�7�7�7�7�78
8888"8(8.848:8@8F8L8R8X8^8d8j8r8x8~8  �0�011"1'1c1�13=3�3�3�3�3�3�3�3�3�3�445J52U2a2|2�2)3�5�5�56#6C6c6�6�6�6	7747J7P7V7\7b7h7n7t7z7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 �  �   L0P0T0X0d0x0|0�0�0�0�0�0�0�01101@1L1P1\1h1t1x1�1�1�1�1�1�1�1�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 444444484X4x4�4�4�4�45�;   �     �7�7�7�7�7�7�78888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�:�:�:�:�:�:H;L;  1�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3�7�7�7�7�7�7�7�7�7�7�7�7�7 �  <   �0�0�0�0l1�1�1�1D2d2�1$2�2�2�:;; ;4;<;L;`;p;|;�;                                                                                                                                                                                                                                                                  